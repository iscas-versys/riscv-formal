`define SYNTHESIS