`ifndef VERILATOR
module testbench;
  reg [4095:0] vcdfile;
  reg clock;
`else
module testbench(input clock, output reg genclock);
  initial genclock = 1;
`endif
  reg genclock = 1;
  reg [31:0] cycle = 0;
  reg [0:0] PI_reset;
  wire [0:0] PI_clock = clock;
  rvfi_testbench UUT (
    .reset(PI_reset),
    .clock(PI_clock)
  );
`ifndef VERILATOR
  initial begin
    if ($value$plusargs("vcd=%s", vcdfile)) begin
      $dumpfile(vcdfile);
      $dumpvars(0, testbench);
    end
    #5 clock = 0;
    while (genclock) begin
      #5 clock = 0;
      #5 clock = 1;
    end
  end
`endif
  initial begin
`ifndef VERILATOR
    #1;
`endif
    UUT.cycle_reg = 8'b00000000;
    UUT.wrapper.core_reset = 1'b1;
    UUT.wrapper.counter = 2'b00;
    UUT.wrapper.uut.core.REG = 1'b0;
    UUT.wrapper.uut.core.REG_1 = 1'b0;
    UUT.wrapper.uut.core.REG_2 = 1'b0;
    UUT.wrapper.uut.core.REG_4 = 1'b1;
    UUT.wrapper.uut.core.REG_5 = 10'b0000001101;
    UUT.wrapper.uut.core.REG_6 = 10'b1111101111;
    UUT.wrapper.uut.core.alu_exe_unit.ALUUnit.r_data_0 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.alu_exe_unit.ALUUnit.r_data_1 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.alu_exe_unit.ALUUnit.r_data_2 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    UUT.wrapper.uut.core.alu_exe_unit.ALUUnit.r_uops_0_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.alu_exe_unit.ALUUnit.r_uops_0_bypassable = 1'b0;
    UUT.wrapper.uut.core.alu_exe_unit.ALUUnit.r_uops_0_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.alu_exe_unit.ALUUnit.r_uops_0_is_amo = 1'b0;
    UUT.wrapper.uut.core.alu_exe_unit.ALUUnit.r_uops_0_pdst = 7'b0000000;
    UUT.wrapper.uut.core.alu_exe_unit.ALUUnit.r_uops_0_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.alu_exe_unit.ALUUnit.r_uops_0_uses_stq = 1'b0;
    UUT.wrapper.uut.core.alu_exe_unit.ALUUnit.r_uops_1_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.alu_exe_unit.ALUUnit.r_uops_1_bypassable = 1'b0;
    UUT.wrapper.uut.core.alu_exe_unit.ALUUnit.r_uops_1_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.alu_exe_unit.ALUUnit.r_uops_1_is_amo = 1'b0;
    UUT.wrapper.uut.core.alu_exe_unit.ALUUnit.r_uops_1_pdst = 7'b0000000;
    UUT.wrapper.uut.core.alu_exe_unit.ALUUnit.r_uops_1_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.alu_exe_unit.ALUUnit.r_uops_1_uses_stq = 1'b0;
    UUT.wrapper.uut.core.alu_exe_unit.ALUUnit.r_uops_2_br_mask = 12'b111111111111;
    UUT.wrapper.uut.core.alu_exe_unit.ALUUnit.r_uops_2_bypassable = 1'b0;
    UUT.wrapper.uut.core.alu_exe_unit.ALUUnit.r_uops_2_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.alu_exe_unit.ALUUnit.r_uops_2_is_amo = 1'b0;
    UUT.wrapper.uut.core.alu_exe_unit.ALUUnit.r_uops_2_pdst = 7'b0000000;
    UUT.wrapper.uut.core.alu_exe_unit.ALUUnit.r_uops_2_rob_idx = 6'b000010;
    UUT.wrapper.uut.core.alu_exe_unit.ALUUnit.r_uops_2_uses_stq = 1'b0;
    UUT.wrapper.uut.core.alu_exe_unit.ALUUnit.r_val_0 = 1'b0;
    UUT.wrapper.uut.core.alu_exe_unit.ALUUnit.r_val_1 = 1'b0;
    UUT.wrapper.uut.core.alu_exe_unit.ALUUnit.r_valids_0 = 1'b0;
    UUT.wrapper.uut.core.alu_exe_unit.ALUUnit.r_valids_1 = 1'b0;
    UUT.wrapper.uut.core.alu_exe_unit.ALUUnit.r_valids_2 = 1'b1;
    UUT.wrapper.uut.core.alu_exe_unit.PipelinedMulUnit.imul.in_pipe_b_dw = 1'b1;
    UUT.wrapper.uut.core.alu_exe_unit.PipelinedMulUnit.imul.in_pipe_b_fn = 5'b11111;
    UUT.wrapper.uut.core.alu_exe_unit.PipelinedMulUnit.imul.in_pipe_b_in1 = 64'b1111111111111111111111111111111111111111111111111111111111111111;
    UUT.wrapper.uut.core.alu_exe_unit.PipelinedMulUnit.imul.in_pipe_b_in2 = 64'b1111111111111111111111111111111111111111111111111111111111111111;
    UUT.wrapper.uut.core.alu_exe_unit.PipelinedMulUnit.imul.in_pipe_v = 1'b0;
    UUT.wrapper.uut.core.alu_exe_unit.PipelinedMulUnit.imul.io_resp_bits_data_pipe_b = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.alu_exe_unit.PipelinedMulUnit.imul.io_resp_bits_data_pipe_pipe_b = 64'b0000000000000000000000000000000000000000000000000000000000010000;
    UUT.wrapper.uut.core.alu_exe_unit.PipelinedMulUnit.imul.io_resp_bits_data_pipe_v = 1'b1;
    UUT.wrapper.uut.core.alu_exe_unit.PipelinedMulUnit.r_uops_0_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.alu_exe_unit.PipelinedMulUnit.r_uops_0_bypassable = 1'b0;
    UUT.wrapper.uut.core.alu_exe_unit.PipelinedMulUnit.r_uops_0_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.alu_exe_unit.PipelinedMulUnit.r_uops_0_is_amo = 1'b0;
    UUT.wrapper.uut.core.alu_exe_unit.PipelinedMulUnit.r_uops_0_pdst = 7'b0000000;
    UUT.wrapper.uut.core.alu_exe_unit.PipelinedMulUnit.r_uops_0_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.alu_exe_unit.PipelinedMulUnit.r_uops_0_uses_stq = 1'b0;
    UUT.wrapper.uut.core.alu_exe_unit.PipelinedMulUnit.r_uops_1_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.alu_exe_unit.PipelinedMulUnit.r_uops_1_bypassable = 1'b0;
    UUT.wrapper.uut.core.alu_exe_unit.PipelinedMulUnit.r_uops_1_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.alu_exe_unit.PipelinedMulUnit.r_uops_1_is_amo = 1'b0;
    UUT.wrapper.uut.core.alu_exe_unit.PipelinedMulUnit.r_uops_1_pdst = 7'b0000000;
    UUT.wrapper.uut.core.alu_exe_unit.PipelinedMulUnit.r_uops_1_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.alu_exe_unit.PipelinedMulUnit.r_uops_1_uses_stq = 1'b0;
    UUT.wrapper.uut.core.alu_exe_unit.PipelinedMulUnit.r_uops_2_br_mask = 12'b111111111111;
    UUT.wrapper.uut.core.alu_exe_unit.PipelinedMulUnit.r_uops_2_bypassable = 1'b0;
    UUT.wrapper.uut.core.alu_exe_unit.PipelinedMulUnit.r_uops_2_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.alu_exe_unit.PipelinedMulUnit.r_uops_2_is_amo = 1'b0;
    UUT.wrapper.uut.core.alu_exe_unit.PipelinedMulUnit.r_uops_2_pdst = 7'b0000000;
    UUT.wrapper.uut.core.alu_exe_unit.PipelinedMulUnit.r_uops_2_rob_idx = 6'b000010;
    UUT.wrapper.uut.core.alu_exe_unit.PipelinedMulUnit.r_uops_2_uses_stq = 1'b0;
    UUT.wrapper.uut.core.alu_exe_unit.PipelinedMulUnit.r_valids_0 = 1'b0;
    UUT.wrapper.uut.core.alu_exe_unit.PipelinedMulUnit.r_valids_1 = 1'b0;
    UUT.wrapper.uut.core.alu_exe_unit.PipelinedMulUnit.r_valids_2 = 1'b1;
    UUT.wrapper.uut.core.alu_exe_unit_1.ALUUnit.r_data_0 = 64'b0000000000000000000000000010000001000000010001000000100000010100;
    UUT.wrapper.uut.core.alu_exe_unit_1.ALUUnit.r_uops_0_br_mask = 12'b111111111111;
    UUT.wrapper.uut.core.alu_exe_unit_1.ALUUnit.r_uops_0_bypassable = 1'b0;
    UUT.wrapper.uut.core.alu_exe_unit_1.ALUUnit.r_uops_0_ctrl_csr_cmd = 3'b010;
    UUT.wrapper.uut.core.alu_exe_unit_1.ALUUnit.r_uops_0_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.alu_exe_unit_1.ALUUnit.r_uops_0_imm_packed = 20'b01111111111111111111;
    UUT.wrapper.uut.core.alu_exe_unit_1.ALUUnit.r_uops_0_is_amo = 1'b0;
    UUT.wrapper.uut.core.alu_exe_unit_1.ALUUnit.r_uops_0_pdst = 7'b0000000;
    UUT.wrapper.uut.core.alu_exe_unit_1.ALUUnit.r_uops_0_rob_idx = 6'b000111;
    UUT.wrapper.uut.core.alu_exe_unit_1.ALUUnit.r_uops_0_uses_stq = 1'b0;
    UUT.wrapper.uut.core.alu_exe_unit_1.ALUUnit.r_valids_0 = 1'b1;
    UUT.wrapper.uut.core.alu_exe_unit_1.DivUnit.div.count = 7'b1111111;
    UUT.wrapper.uut.core.alu_exe_unit_1.DivUnit.div.divisor = 65'b00000000001111111111111111111111111111111111111111111110000000001;
    UUT.wrapper.uut.core.alu_exe_unit_1.DivUnit.div.isHi = 1'b1;
    UUT.wrapper.uut.core.alu_exe_unit_1.DivUnit.div.neg_out = 1'b0;
    UUT.wrapper.uut.core.alu_exe_unit_1.DivUnit.div.remainder = 130'b0000000010000000000000000000000000000000000000000000000000000001010000000010000000000000000000000000000000000000000000000000000010;
    UUT.wrapper.uut.core.alu_exe_unit_1.DivUnit.div.req_dw = 1'b0;
    UUT.wrapper.uut.core.alu_exe_unit_1.DivUnit.div.resHi = 1'b0;
    UUT.wrapper.uut.core.alu_exe_unit_1.DivUnit.div.state = 3'b010;
    UUT.wrapper.uut.core.alu_exe_unit_1.DivUnit.r_uop_br_mask = 12'b111111111111;
    UUT.wrapper.uut.core.alu_exe_unit_1.DivUnit.r_uop_bypassable = 1'b0;
    UUT.wrapper.uut.core.alu_exe_unit_1.DivUnit.r_uop_dst_rtype = 2'b11;
    UUT.wrapper.uut.core.alu_exe_unit_1.DivUnit.r_uop_is_amo = 1'b0;
    UUT.wrapper.uut.core.alu_exe_unit_1.DivUnit.r_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.core.alu_exe_unit_1.DivUnit.r_uop_rob_idx = 6'b000011;
    UUT.wrapper.uut.core.alu_exe_unit_1.DivUnit.r_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.core.alu_exe_unit_io_req_bits_kill_REG = 1'b0;
    UUT.wrapper.uut.core.alu_exe_unit_io_req_bits_kill_REG_1 = 1'b0;
    UUT.wrapper.uut.core.b2_cfi_type = 3'b011;
    UUT.wrapper.uut.core.b2_jalr_target = 40'b0011111111111111111101010111001001111000;
    UUT.wrapper.uut.core.b2_jalr_target_REG = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.b2_mispredict = 1'b0;
    UUT.wrapper.uut.core.b2_pc_sel = 2'b11;
    UUT.wrapper.uut.core.b2_taken = 1'b1;
    UUT.wrapper.uut.core.b2_target_offset = 64'b0000000000000000000000000000000000000000000000000000000000000111;
    UUT.wrapper.uut.core.b2_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.b2_uop_br_tag = 4'b0000;
    UUT.wrapper.uut.core.b2_uop_edge_inst = 1'b0;
    UUT.wrapper.uut.core.b2_uop_ftq_idx = 3'b111;
    UUT.wrapper.uut.core.b2_uop_is_rvc = 1'b1;
    UUT.wrapper.uut.core.b2_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.core.b2_uop_pc_lob = 6'b000001;
    UUT.wrapper.uut.core.b2_uop_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.b2_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.core.brinfos_0_cfi_type = 3'b000;
    UUT.wrapper.uut.core.brinfos_0_mispredict = 1'b0;
    UUT.wrapper.uut.core.brinfos_0_pc_sel = 2'b00;
    UUT.wrapper.uut.core.brinfos_0_taken = 1'b0;
    UUT.wrapper.uut.core.brinfos_0_target_offset = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.brinfos_0_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.brinfos_0_uop_br_tag = 4'b1000;
    UUT.wrapper.uut.core.brinfos_0_uop_edge_inst = 1'b0;
    UUT.wrapper.uut.core.brinfos_0_uop_ftq_idx = 3'b000;
    UUT.wrapper.uut.core.brinfos_0_uop_is_rvc = 1'b0;
    UUT.wrapper.uut.core.brinfos_0_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.core.brinfos_0_uop_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.brinfos_0_uop_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.brinfos_0_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.core.brinfos_0_valid = 1'b1;
    UUT.wrapper.uut.core.brinfos_1_cfi_type = 3'b000;
    UUT.wrapper.uut.core.brinfos_1_mispredict = 1'b0;
    UUT.wrapper.uut.core.brinfos_1_pc_sel = 2'b00;
    UUT.wrapper.uut.core.brinfos_1_taken = 1'b0;
    UUT.wrapper.uut.core.brinfos_1_target_offset = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.brinfos_1_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.brinfos_1_uop_br_tag = 4'b1001;
    UUT.wrapper.uut.core.brinfos_1_uop_edge_inst = 1'b0;
    UUT.wrapper.uut.core.brinfos_1_uop_ftq_idx = 3'b000;
    UUT.wrapper.uut.core.brinfos_1_uop_is_rvc = 1'b0;
    UUT.wrapper.uut.core.brinfos_1_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.core.brinfos_1_uop_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.brinfos_1_uop_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.brinfos_1_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.core.brinfos_1_valid = 1'b1;
    UUT.wrapper.uut.core.csr.io_status_cease_r = 1'b0;
    UUT.wrapper.uut.core.csr.large_ = 58'b1111111111111111111111110000000000000110000000000000111111;
    UUT.wrapper.uut.core.csr.large_1 = 58'b1111111111111111111111111111111111111111111111111111111111;
    UUT.wrapper.uut.core.csr.large_2 = 34'b1111111111111111110111111110000000;
    UUT.wrapper.uut.core.csr.large_3 = 34'b1111111111111111111111111111111111;
    UUT.wrapper.uut.core.csr.large_4 = 34'b0011111111111111111111111111111111;
    UUT.wrapper.uut.core.csr.large_5 = 34'b1111111111011110111111111111000000;
    UUT.wrapper.uut.core.csr.large_6 = 34'b1111010111110111111111111110000000;
    UUT.wrapper.uut.core.csr.large_7 = 34'b1111111101101111110111011110000000;
    UUT.wrapper.uut.core.csr.reg_custom_0 = 64'b0100000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.csr.reg_hpmevent_0 = 64'b1111111111111111111111111111111111111111111111111111010111111101;
    UUT.wrapper.uut.core.csr.reg_hpmevent_1 = 64'b1111111111111111111111111111111111111111111111111111010111111110;
    UUT.wrapper.uut.core.csr.reg_hpmevent_2 = 64'b1111111111111111111111111111111111111111111111111111010111111111;
    UUT.wrapper.uut.core.csr.reg_hpmevent_3 = 64'b1111111111111111111111111111111111111111111111111111010111111111;
    UUT.wrapper.uut.core.csr.reg_hpmevent_4 = 64'b1111111111111111111111111111111111111111111111111111010111111111;
    UUT.wrapper.uut.core.csr.reg_hpmevent_5 = 64'b1111111111111111111111111111111111111111111111111111010111111110;
    UUT.wrapper.uut.core.csr.reg_mcause = 64'b1111111111111111111111111111111111111111111111111111111111111111;
    UUT.wrapper.uut.core.csr.reg_mcounteren = 32'b11111111111111111111111000000000;
    UUT.wrapper.uut.core.csr.reg_mcountinhibit = 9'b111001111;
    UUT.wrapper.uut.core.csr.reg_medeleg = 64'b1111111111111111111111111111111111111111111111110100111010100010;
    UUT.wrapper.uut.core.csr.reg_menvcfg_fiom = 1'b1;
    UUT.wrapper.uut.core.csr.reg_mepc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.csr.reg_mideleg = 64'b0000000000000000000000000000000000000000000000000000001000100010;
    UUT.wrapper.uut.core.csr.reg_mie = 64'b0000000000000000000000000000000000000000000000000000001000101010;
    UUT.wrapper.uut.core.csr.reg_mip_seip = 1'b1;
    UUT.wrapper.uut.core.csr.reg_mip_ssip = 1'b1;
    UUT.wrapper.uut.core.csr.reg_mip_stip = 1'b1;
    UUT.wrapper.uut.core.csr.reg_mscratch = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.csr.reg_mstatus_fs = 2'b11;
    UUT.wrapper.uut.core.csr.reg_mstatus_mie = 1'b0;
    UUT.wrapper.uut.core.csr.reg_mstatus_mpie = 1'b0;
    UUT.wrapper.uut.core.csr.reg_mstatus_mpp = 2'b01;
    UUT.wrapper.uut.core.csr.reg_mstatus_mprv = 1'b1;
    UUT.wrapper.uut.core.csr.reg_mstatus_mxr = 1'b1;
    UUT.wrapper.uut.core.csr.reg_mstatus_prv = 2'b11;
    UUT.wrapper.uut.core.csr.reg_mstatus_sie = 1'b1;
    UUT.wrapper.uut.core.csr.reg_mstatus_spie = 1'b1;
    UUT.wrapper.uut.core.csr.reg_mstatus_spp = 1'b1;
    UUT.wrapper.uut.core.csr.reg_mstatus_sum = 1'b0;
    UUT.wrapper.uut.core.csr.reg_mstatus_tsr = 1'b0;
    UUT.wrapper.uut.core.csr.reg_mstatus_tvm = 1'b0;
    UUT.wrapper.uut.core.csr.reg_mstatus_tw = 1'b0;
    UUT.wrapper.uut.core.csr.reg_mtval = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.csr.reg_mtvec = 32'b00000000000000000000000011111011;
    UUT.wrapper.uut.core.csr.reg_satp_mode = 4'b1111;
    UUT.wrapper.uut.core.csr.reg_satp_ppn = 44'b11111111111111111111111100000000000000000000;
    UUT.wrapper.uut.core.csr.reg_scause = 64'b0000000000000000000000000000000000000000000000000000000011100000;
    UUT.wrapper.uut.core.csr.reg_scounteren = 32'b11111111111111111111111000000000;
    UUT.wrapper.uut.core.csr.reg_senvcfg_fiom = 1'b1;
    UUT.wrapper.uut.core.csr.reg_sepc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.csr.reg_singleStepped = 1'b0;
    UUT.wrapper.uut.core.csr.reg_sscratch = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.csr.reg_stval = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.csr.reg_stvec = 39'b000000000000000000000000000000000000011;
    UUT.wrapper.uut.core.csr.reg_wfi = 1'b0;
    UUT.wrapper.uut.core.csr.small_ = 6'b001001;
    UUT.wrapper.uut.core.csr.small_1 = 6'b111111;
    UUT.wrapper.uut.core.csr.small_2 = 6'b111111;
    UUT.wrapper.uut.core.csr.small_3 = 6'b111111;
    UUT.wrapper.uut.core.csr.small_4 = 6'b111111;
    UUT.wrapper.uut.core.csr.small_5 = 6'b111111;
    UUT.wrapper.uut.core.csr.small_6 = 6'b111111;
    UUT.wrapper.uut.core.csr.small_7 = 6'b011111;
    UUT.wrapper.uut.core.csr_io_cause_REG = 64'b1000000000000000000000000000000000000000000000000000000011110111;
    UUT.wrapper.uut.core.csr_io_counters_0_inc_REG = 1'b1;
    UUT.wrapper.uut.core.csr_io_counters_1_inc_REG = 1'b1;
    UUT.wrapper.uut.core.csr_io_counters_2_inc_REG = 1'b1;
    UUT.wrapper.uut.core.csr_io_counters_3_inc_REG = 1'b1;
    UUT.wrapper.uut.core.csr_io_counters_4_inc_REG = 1'b1;
    UUT.wrapper.uut.core.csr_io_counters_5_inc_REG = 1'b1;
    UUT.wrapper.uut.core.csr_io_exception_REG = 1'b0;
    UUT.wrapper.uut.core.csr_io_pc_REG = 6'b000001;
    UUT.wrapper.uut.core.csr_io_pc_REG_1 = 1'b0;
    UUT.wrapper.uut.core.csr_io_retire_REG = 2'b00;
    UUT.wrapper.uut.core.csr_io_tval_REG = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_0_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_0_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_0_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_0_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_10_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_10_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_10_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_10_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_11_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_11_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_11_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_11_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_12_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_12_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_12_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_12_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_13_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_13_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_13_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_13_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_14_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_14_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_14_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_14_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_15_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_15_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_15_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_15_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_16_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_16_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_16_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_16_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_17_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_17_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_17_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_17_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_18_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_18_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_18_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_18_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_19_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_19_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_19_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_19_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_1_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_1_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_1_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_1_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_20_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_20_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_20_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_20_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_21_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_21_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_21_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_21_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_22_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_22_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_22_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_22_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_23_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_23_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_23_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_23_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_24_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_24_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_24_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_24_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_25_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_25_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_25_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_25_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_26_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_26_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_26_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_26_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_27_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_27_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_27_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_27_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_28_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_28_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_28_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_28_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_29_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_29_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_29_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_29_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_2_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_2_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_2_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_2_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_30_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_30_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_30_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_30_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_31_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_31_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_31_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_31_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_32_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_32_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_32_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_32_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_33_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_33_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_33_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_33_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_34_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_34_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_34_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_34_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_35_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_35_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_35_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_35_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_36_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_36_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_36_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_36_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_37_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_37_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_37_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_37_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_38_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_38_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_38_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_38_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_39_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_39_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_39_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_39_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_3_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_3_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_3_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_3_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_40_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_40_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_40_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_40_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_41_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_41_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_41_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_41_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_42_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_42_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_42_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_42_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_43_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_43_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_43_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_43_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_44_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_44_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_44_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_44_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_45_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_45_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_45_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_45_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_46_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_46_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_46_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_46_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_47_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_47_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_47_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_47_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_48_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_48_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_48_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_48_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_49_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_49_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_49_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_49_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_4_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_4_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_4_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_4_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_50_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_50_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_50_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_50_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_51_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_51_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_51_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_51_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_52_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_52_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_52_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_52_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_53_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_53_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_53_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_53_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_54_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_54_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_54_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_54_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_55_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_55_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_55_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_55_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_56_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_56_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_56_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_56_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_57_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_57_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_57_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_57_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_58_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_58_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_58_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_58_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_59_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_59_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_59_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_59_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_5_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_5_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_5_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_5_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_60_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_60_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_60_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_60_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_61_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_61_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_61_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_61_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_62_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_62_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_62_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_62_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_63_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_63_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_63_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_63_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_6_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_6_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_6_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_6_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_7_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_7_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_7_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_7_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_8_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_8_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_8_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_8_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_9_cfi_type = 3'b000;
    UUT.wrapper.uut.core.debug_br_res_9_jalr_target = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_9_target_offset = 21'b000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_9_valid = 1'b0;
    UUT.wrapper.uut.core.debug_br_res_jalr_target_REG = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.debug_br_res_jalr_target_REG_1 = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.dec_brmask_logic.branch_mask = 12'b000000000000;
    UUT.wrapper.uut.core.dec_brmask_logic_io_flush_pipeline_REG = 1'b0;
    UUT.wrapper.uut.core.dec_finished_mask = 2'b00;
    UUT.wrapper.uut.core.flush_pc_REG = 6'b111100;
    UUT.wrapper.uut.core.flush_pc_REG_1 = 1'b0;
    UUT.wrapper.uut.core.flush_pc_next_REG = 1'b0;
    UUT.wrapper.uut.core.flush_typ = 3'b011;
    UUT.wrapper.uut.core.int_issue_unit.io_dis_uops_0_ready_REG = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.io_dis_uops_1_ready_REG = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_0.p1 = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_0.p1_poisoned = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_0.p2 = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_0.p2_poisoned = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_0.p3 = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_0.ppred = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_0.slot_uop_br_mask = 12'b111111111111;
    UUT.wrapper.uut.core.int_issue_unit.slots_0.slot_uop_br_tag = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_0.slot_uop_bypassable = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_0.slot_uop_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_0.slot_uop_edge_inst = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_0.slot_uop_ftq_idx = 3'b000;
    UUT.wrapper.uut.core.int_issue_unit.slots_0.slot_uop_fu_code = 10'b1111000101;
    UUT.wrapper.uut.core.int_issue_unit.slots_0.slot_uop_imm_packed = 20'b00000000000000000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_0.slot_uop_is_amo = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_0.slot_uop_is_br = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_0.slot_uop_is_jal = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_0.slot_uop_is_jalr = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_0.slot_uop_is_rvc = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_0.slot_uop_is_sfb = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_0.slot_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_0.slot_uop_ldst_val = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_0.slot_uop_lrs1_rtype = 2'b11;
    UUT.wrapper.uut.core.int_issue_unit.slots_0.slot_uop_lrs2_rtype = 2'b11;
    UUT.wrapper.uut.core.int_issue_unit.slots_0.slot_uop_mem_cmd = 5'b00000;
    UUT.wrapper.uut.core.int_issue_unit.slots_0.slot_uop_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_0.slot_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_0.slot_uop_prs1 = 7'b1111111;
    UUT.wrapper.uut.core.int_issue_unit.slots_0.slot_uop_prs2 = 7'b1111111;
    UUT.wrapper.uut.core.int_issue_unit.slots_0.slot_uop_prs3 = 7'b1111111;
    UUT.wrapper.uut.core.int_issue_unit.slots_0.slot_uop_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_0.slot_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_0.slot_uop_taken = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_0.slot_uop_uopc = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_0.slot_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_0.state = 2'b10;
    UUT.wrapper.uut.core.int_issue_unit.slots_1.p1 = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_1.p1_poisoned = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_1.p2 = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_1.p2_poisoned = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_1.p3 = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_1.ppred = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_1.slot_uop_br_mask = 12'b111111111111;
    UUT.wrapper.uut.core.int_issue_unit.slots_1.slot_uop_br_tag = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_1.slot_uop_bypassable = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_1.slot_uop_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_1.slot_uop_edge_inst = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_1.slot_uop_ftq_idx = 3'b000;
    UUT.wrapper.uut.core.int_issue_unit.slots_1.slot_uop_fu_code = 10'b1111000100;
    UUT.wrapper.uut.core.int_issue_unit.slots_1.slot_uop_imm_packed = 20'b00000000000000000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_1.slot_uop_is_amo = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_1.slot_uop_is_br = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_1.slot_uop_is_jal = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_1.slot_uop_is_jalr = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_1.slot_uop_is_rvc = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_1.slot_uop_is_sfb = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_1.slot_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_1.slot_uop_ldst_val = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_1.slot_uop_lrs1_rtype = 2'b11;
    UUT.wrapper.uut.core.int_issue_unit.slots_1.slot_uop_lrs2_rtype = 2'b11;
    UUT.wrapper.uut.core.int_issue_unit.slots_1.slot_uop_mem_cmd = 5'b00000;
    UUT.wrapper.uut.core.int_issue_unit.slots_1.slot_uop_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_1.slot_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_1.slot_uop_prs1 = 7'b1111111;
    UUT.wrapper.uut.core.int_issue_unit.slots_1.slot_uop_prs2 = 7'b1111111;
    UUT.wrapper.uut.core.int_issue_unit.slots_1.slot_uop_prs3 = 7'b1111111;
    UUT.wrapper.uut.core.int_issue_unit.slots_1.slot_uop_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_1.slot_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_1.slot_uop_taken = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_1.slot_uop_uopc = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_1.slot_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_1.state = 2'b10;
    UUT.wrapper.uut.core.int_issue_unit.slots_10.p1 = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_10.p1_poisoned = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_10.p2 = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_10.p2_poisoned = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_10.p3 = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_10.ppred = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_10.slot_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_10.slot_uop_br_tag = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_10.slot_uop_bypassable = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_10.slot_uop_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_10.slot_uop_edge_inst = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_10.slot_uop_ftq_idx = 3'b000;
    UUT.wrapper.uut.core.int_issue_unit.slots_10.slot_uop_fu_code = 10'b0000000001;
    UUT.wrapper.uut.core.int_issue_unit.slots_10.slot_uop_imm_packed = 20'b00000000000000000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_10.slot_uop_is_amo = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_10.slot_uop_is_br = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_10.slot_uop_is_jal = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_10.slot_uop_is_jalr = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_10.slot_uop_is_rvc = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_10.slot_uop_is_sfb = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_10.slot_uop_ldq_idx = 4'b1111;
    UUT.wrapper.uut.core.int_issue_unit.slots_10.slot_uop_ldst_val = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_10.slot_uop_lrs1_rtype = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_10.slot_uop_lrs2_rtype = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_10.slot_uop_mem_cmd = 5'b00000;
    UUT.wrapper.uut.core.int_issue_unit.slots_10.slot_uop_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_10.slot_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_10.slot_uop_prs1 = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_10.slot_uop_prs2 = 7'b0000011;
    UUT.wrapper.uut.core.int_issue_unit.slots_10.slot_uop_prs3 = 7'b0000010;
    UUT.wrapper.uut.core.int_issue_unit.slots_10.slot_uop_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_10.slot_uop_stq_idx = 4'b1111;
    UUT.wrapper.uut.core.int_issue_unit.slots_10.slot_uop_taken = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_10.slot_uop_uopc = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_10.slot_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_10.state = 2'b01;
    UUT.wrapper.uut.core.int_issue_unit.slots_11.p1 = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_11.p1_poisoned = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_11.p2 = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_11.p2_poisoned = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_11.p3 = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_11.ppred = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_11.slot_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_11.slot_uop_br_tag = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_11.slot_uop_bypassable = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_11.slot_uop_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_11.slot_uop_edge_inst = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_11.slot_uop_ftq_idx = 3'b001;
    UUT.wrapper.uut.core.int_issue_unit.slots_11.slot_uop_fu_code = 10'b0000011011;
    UUT.wrapper.uut.core.int_issue_unit.slots_11.slot_uop_imm_packed = 20'b00000010000000000100;
    UUT.wrapper.uut.core.int_issue_unit.slots_11.slot_uop_is_amo = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_11.slot_uop_is_br = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_11.slot_uop_is_jal = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_11.slot_uop_is_jalr = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_11.slot_uop_is_rvc = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_11.slot_uop_is_sfb = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_11.slot_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_11.slot_uop_ldst_val = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_11.slot_uop_lrs1_rtype = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_11.slot_uop_lrs2_rtype = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_11.slot_uop_mem_cmd = 5'b00000;
    UUT.wrapper.uut.core.int_issue_unit.slots_11.slot_uop_pc_lob = 6'b000100;
    UUT.wrapper.uut.core.int_issue_unit.slots_11.slot_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_11.slot_uop_prs1 = 7'b0000010;
    UUT.wrapper.uut.core.int_issue_unit.slots_11.slot_uop_prs2 = 7'b0000010;
    UUT.wrapper.uut.core.int_issue_unit.slots_11.slot_uop_prs3 = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_11.slot_uop_rob_idx = 6'b000010;
    UUT.wrapper.uut.core.int_issue_unit.slots_11.slot_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_11.slot_uop_taken = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_11.slot_uop_uopc = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_11.slot_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_11.state = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_12.p1 = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_12.p1_poisoned = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_12.p2 = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_12.p2_poisoned = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_12.p3 = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_12.ppred = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_12.slot_uop_br_mask = 12'b000000000001;
    UUT.wrapper.uut.core.int_issue_unit.slots_12.slot_uop_br_tag = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_12.slot_uop_bypassable = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_12.slot_uop_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_12.slot_uop_edge_inst = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_12.slot_uop_ftq_idx = 3'b000;
    UUT.wrapper.uut.core.int_issue_unit.slots_12.slot_uop_fu_code = 10'b0000000001;
    UUT.wrapper.uut.core.int_issue_unit.slots_12.slot_uop_imm_packed = 20'b00000010000000110110;
    UUT.wrapper.uut.core.int_issue_unit.slots_12.slot_uop_is_amo = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_12.slot_uop_is_br = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_12.slot_uop_is_jal = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_12.slot_uop_is_jalr = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_12.slot_uop_is_rvc = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_12.slot_uop_is_sfb = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_12.slot_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_12.slot_uop_ldst_val = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_12.slot_uop_lrs1_rtype = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_12.slot_uop_lrs2_rtype = 2'b01;
    UUT.wrapper.uut.core.int_issue_unit.slots_12.slot_uop_mem_cmd = 5'b00000;
    UUT.wrapper.uut.core.int_issue_unit.slots_12.slot_uop_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_12.slot_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_12.slot_uop_prs1 = 7'b0000111;
    UUT.wrapper.uut.core.int_issue_unit.slots_12.slot_uop_prs2 = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_12.slot_uop_prs3 = 7'b0000010;
    UUT.wrapper.uut.core.int_issue_unit.slots_12.slot_uop_rob_idx = 6'b000010;
    UUT.wrapper.uut.core.int_issue_unit.slots_12.slot_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_12.slot_uop_taken = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_12.slot_uop_uopc = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_12.slot_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_12.state = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_13.p1 = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_13.p1_poisoned = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_13.p2 = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_13.p2_poisoned = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_13.p3 = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_13.ppred = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_13.slot_uop_br_mask = 12'b000000000010;
    UUT.wrapper.uut.core.int_issue_unit.slots_13.slot_uop_br_tag = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_13.slot_uop_bypassable = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_13.slot_uop_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_13.slot_uop_edge_inst = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_13.slot_uop_ftq_idx = 3'b010;
    UUT.wrapper.uut.core.int_issue_unit.slots_13.slot_uop_fu_code = 10'b0000010000;
    UUT.wrapper.uut.core.int_issue_unit.slots_13.slot_uop_imm_packed = 20'b00000010000000000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_13.slot_uop_is_amo = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_13.slot_uop_is_br = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_13.slot_uop_is_jal = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_13.slot_uop_is_jalr = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_13.slot_uop_is_rvc = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_13.slot_uop_is_sfb = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_13.slot_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_13.slot_uop_ldst_val = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_13.slot_uop_lrs1_rtype = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_13.slot_uop_lrs2_rtype = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_13.slot_uop_mem_cmd = 5'b00000;
    UUT.wrapper.uut.core.int_issue_unit.slots_13.slot_uop_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_13.slot_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_13.slot_uop_prs1 = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_13.slot_uop_prs2 = 7'b1000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_13.slot_uop_prs3 = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_13.slot_uop_rob_idx = 6'b000011;
    UUT.wrapper.uut.core.int_issue_unit.slots_13.slot_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_13.slot_uop_taken = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_13.slot_uop_uopc = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_13.slot_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_13.state = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_14.p1 = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_14.p1_poisoned = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_14.p2 = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_14.p2_poisoned = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_14.p3 = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_14.ppred = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_14.slot_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_14.slot_uop_br_tag = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_14.slot_uop_bypassable = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_14.slot_uop_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_14.slot_uop_edge_inst = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_14.slot_uop_ftq_idx = 3'b000;
    UUT.wrapper.uut.core.int_issue_unit.slots_14.slot_uop_fu_code = 10'b0000000001;
    UUT.wrapper.uut.core.int_issue_unit.slots_14.slot_uop_imm_packed = 20'b00000010001111110110;
    UUT.wrapper.uut.core.int_issue_unit.slots_14.slot_uop_is_amo = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_14.slot_uop_is_br = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_14.slot_uop_is_jal = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_14.slot_uop_is_jalr = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_14.slot_uop_is_rvc = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_14.slot_uop_is_sfb = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_14.slot_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_14.slot_uop_ldst_val = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_14.slot_uop_lrs1_rtype = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_14.slot_uop_lrs2_rtype = 2'b11;
    UUT.wrapper.uut.core.int_issue_unit.slots_14.slot_uop_mem_cmd = 5'b00000;
    UUT.wrapper.uut.core.int_issue_unit.slots_14.slot_uop_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_14.slot_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_14.slot_uop_prs1 = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_14.slot_uop_prs2 = 7'b0000001;
    UUT.wrapper.uut.core.int_issue_unit.slots_14.slot_uop_prs3 = 7'b0000011;
    UUT.wrapper.uut.core.int_issue_unit.slots_14.slot_uop_rob_idx = 6'b000010;
    UUT.wrapper.uut.core.int_issue_unit.slots_14.slot_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_14.slot_uop_taken = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_14.slot_uop_uopc = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_14.slot_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_14.state = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_15.p1 = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_15.p1_poisoned = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_15.p2 = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_15.p2_poisoned = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_15.p3 = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_15.ppred = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_15.slot_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_15.slot_uop_br_tag = 4'b0010;
    UUT.wrapper.uut.core.int_issue_unit.slots_15.slot_uop_bypassable = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_15.slot_uop_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_15.slot_uop_edge_inst = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_15.slot_uop_ftq_idx = 3'b010;
    UUT.wrapper.uut.core.int_issue_unit.slots_15.slot_uop_fu_code = 10'b0000000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_15.slot_uop_imm_packed = 20'b00000000000000000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_15.slot_uop_is_amo = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_15.slot_uop_is_br = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_15.slot_uop_is_jal = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_15.slot_uop_is_jalr = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_15.slot_uop_is_rvc = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_15.slot_uop_is_sfb = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_15.slot_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_15.slot_uop_ldst_val = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_15.slot_uop_lrs1_rtype = 2'b01;
    UUT.wrapper.uut.core.int_issue_unit.slots_15.slot_uop_lrs2_rtype = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_15.slot_uop_mem_cmd = 5'b00000;
    UUT.wrapper.uut.core.int_issue_unit.slots_15.slot_uop_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_15.slot_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_15.slot_uop_prs1 = 7'b0001000;
    UUT.wrapper.uut.core.int_issue_unit.slots_15.slot_uop_prs2 = 7'b1000010;
    UUT.wrapper.uut.core.int_issue_unit.slots_15.slot_uop_prs3 = 7'b0000100;
    UUT.wrapper.uut.core.int_issue_unit.slots_15.slot_uop_rob_idx = 6'b000011;
    UUT.wrapper.uut.core.int_issue_unit.slots_15.slot_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_15.slot_uop_taken = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_15.slot_uop_uopc = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_15.slot_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_15.state = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_16.p1 = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_16.p1_poisoned = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_16.p2 = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_16.p2_poisoned = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_16.p3 = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_16.ppred = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_16.slot_uop_br_mask = 12'b001100000001;
    UUT.wrapper.uut.core.int_issue_unit.slots_16.slot_uop_br_tag = 4'b0001;
    UUT.wrapper.uut.core.int_issue_unit.slots_16.slot_uop_bypassable = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_16.slot_uop_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_16.slot_uop_edge_inst = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_16.slot_uop_ftq_idx = 3'b000;
    UUT.wrapper.uut.core.int_issue_unit.slots_16.slot_uop_fu_code = 10'b0000000001;
    UUT.wrapper.uut.core.int_issue_unit.slots_16.slot_uop_imm_packed = 20'b00000010000000110010;
    UUT.wrapper.uut.core.int_issue_unit.slots_16.slot_uop_is_amo = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_16.slot_uop_is_br = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_16.slot_uop_is_jal = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_16.slot_uop_is_jalr = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_16.slot_uop_is_rvc = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_16.slot_uop_is_sfb = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_16.slot_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_16.slot_uop_ldst_val = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_16.slot_uop_lrs1_rtype = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_16.slot_uop_lrs2_rtype = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_16.slot_uop_mem_cmd = 5'b00000;
    UUT.wrapper.uut.core.int_issue_unit.slots_16.slot_uop_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_16.slot_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_16.slot_uop_prs1 = 7'b0000001;
    UUT.wrapper.uut.core.int_issue_unit.slots_16.slot_uop_prs2 = 7'b0000001;
    UUT.wrapper.uut.core.int_issue_unit.slots_16.slot_uop_prs3 = 7'b0000001;
    UUT.wrapper.uut.core.int_issue_unit.slots_16.slot_uop_rob_idx = 6'b000010;
    UUT.wrapper.uut.core.int_issue_unit.slots_16.slot_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_16.slot_uop_taken = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_16.slot_uop_uopc = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_16.slot_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_16.state = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_17.p1 = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_17.p1_poisoned = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_17.p2 = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_17.p2_poisoned = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_17.p3 = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_17.ppred = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_17.slot_uop_br_mask = 12'b001100000001;
    UUT.wrapper.uut.core.int_issue_unit.slots_17.slot_uop_br_tag = 4'b0001;
    UUT.wrapper.uut.core.int_issue_unit.slots_17.slot_uop_bypassable = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_17.slot_uop_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_17.slot_uop_edge_inst = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_17.slot_uop_ftq_idx = 3'b001;
    UUT.wrapper.uut.core.int_issue_unit.slots_17.slot_uop_fu_code = 10'b0000001010;
    UUT.wrapper.uut.core.int_issue_unit.slots_17.slot_uop_imm_packed = 20'b00000000100000000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_17.slot_uop_is_amo = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_17.slot_uop_is_br = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_17.slot_uop_is_jal = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_17.slot_uop_is_jalr = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_17.slot_uop_is_rvc = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_17.slot_uop_is_sfb = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_17.slot_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_17.slot_uop_ldst_val = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_17.slot_uop_lrs1_rtype = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_17.slot_uop_lrs2_rtype = 2'b01;
    UUT.wrapper.uut.core.int_issue_unit.slots_17.slot_uop_mem_cmd = 5'b00000;
    UUT.wrapper.uut.core.int_issue_unit.slots_17.slot_uop_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_17.slot_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_17.slot_uop_prs1 = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_17.slot_uop_prs2 = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_17.slot_uop_prs3 = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_17.slot_uop_rob_idx = 6'b000001;
    UUT.wrapper.uut.core.int_issue_unit.slots_17.slot_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_17.slot_uop_taken = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_17.slot_uop_uopc = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_17.slot_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_17.state = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_18.p1 = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_18.p1_poisoned = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_18.p2 = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_18.p2_poisoned = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_18.p3 = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_18.ppred = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_18.slot_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_18.slot_uop_br_tag = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_18.slot_uop_bypassable = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_18.slot_uop_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_18.slot_uop_edge_inst = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_18.slot_uop_ftq_idx = 3'b000;
    UUT.wrapper.uut.core.int_issue_unit.slots_18.slot_uop_fu_code = 10'b0000111011;
    UUT.wrapper.uut.core.int_issue_unit.slots_18.slot_uop_imm_packed = 20'b00000000000000000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_18.slot_uop_is_amo = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_18.slot_uop_is_br = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_18.slot_uop_is_jal = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_18.slot_uop_is_jalr = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_18.slot_uop_is_rvc = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_18.slot_uop_is_sfb = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_18.slot_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_18.slot_uop_ldst_val = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_18.slot_uop_lrs1_rtype = 2'b01;
    UUT.wrapper.uut.core.int_issue_unit.slots_18.slot_uop_lrs2_rtype = 2'b01;
    UUT.wrapper.uut.core.int_issue_unit.slots_18.slot_uop_mem_cmd = 5'b00000;
    UUT.wrapper.uut.core.int_issue_unit.slots_18.slot_uop_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_18.slot_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_18.slot_uop_prs1 = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_18.slot_uop_prs2 = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_18.slot_uop_prs3 = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_18.slot_uop_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_18.slot_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_18.slot_uop_taken = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_18.slot_uop_uopc = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_18.slot_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_18.state = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_19.p1 = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_19.p1_poisoned = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_19.p2 = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_19.p2_poisoned = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_19.p3 = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_19.ppred = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_19.slot_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_19.slot_uop_br_tag = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_19.slot_uop_bypassable = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_19.slot_uop_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_19.slot_uop_edge_inst = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_19.slot_uop_ftq_idx = 3'b000;
    UUT.wrapper.uut.core.int_issue_unit.slots_19.slot_uop_fu_code = 10'b0000111011;
    UUT.wrapper.uut.core.int_issue_unit.slots_19.slot_uop_imm_packed = 20'b00000000000000000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_19.slot_uop_is_amo = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_19.slot_uop_is_br = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_19.slot_uop_is_jal = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_19.slot_uop_is_jalr = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_19.slot_uop_is_rvc = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_19.slot_uop_is_sfb = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_19.slot_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_19.slot_uop_ldst_val = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_19.slot_uop_lrs1_rtype = 2'b01;
    UUT.wrapper.uut.core.int_issue_unit.slots_19.slot_uop_lrs2_rtype = 2'b01;
    UUT.wrapper.uut.core.int_issue_unit.slots_19.slot_uop_mem_cmd = 5'b00000;
    UUT.wrapper.uut.core.int_issue_unit.slots_19.slot_uop_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_19.slot_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_19.slot_uop_prs1 = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_19.slot_uop_prs2 = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_19.slot_uop_prs3 = 7'b1111111;
    UUT.wrapper.uut.core.int_issue_unit.slots_19.slot_uop_rob_idx = 6'b111111;
    UUT.wrapper.uut.core.int_issue_unit.slots_19.slot_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_19.slot_uop_taken = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_19.slot_uop_uopc = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_19.slot_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_19.state = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_2.p1 = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_2.p1_poisoned = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_2.p2 = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_2.p2_poisoned = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_2.p3 = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_2.ppred = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_2.slot_uop_br_mask = 12'b111111111111;
    UUT.wrapper.uut.core.int_issue_unit.slots_2.slot_uop_br_tag = 4'b1111;
    UUT.wrapper.uut.core.int_issue_unit.slots_2.slot_uop_bypassable = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_2.slot_uop_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_2.slot_uop_edge_inst = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_2.slot_uop_ftq_idx = 3'b111;
    UUT.wrapper.uut.core.int_issue_unit.slots_2.slot_uop_fu_code = 10'b1111000100;
    UUT.wrapper.uut.core.int_issue_unit.slots_2.slot_uop_imm_packed = 20'b11111111111111111111;
    UUT.wrapper.uut.core.int_issue_unit.slots_2.slot_uop_is_amo = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_2.slot_uop_is_br = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_2.slot_uop_is_jal = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_2.slot_uop_is_jalr = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_2.slot_uop_is_rvc = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_2.slot_uop_is_sfb = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_2.slot_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_2.slot_uop_ldst_val = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_2.slot_uop_lrs1_rtype = 2'b11;
    UUT.wrapper.uut.core.int_issue_unit.slots_2.slot_uop_lrs2_rtype = 2'b11;
    UUT.wrapper.uut.core.int_issue_unit.slots_2.slot_uop_mem_cmd = 5'b11111;
    UUT.wrapper.uut.core.int_issue_unit.slots_2.slot_uop_pc_lob = 6'b111111;
    UUT.wrapper.uut.core.int_issue_unit.slots_2.slot_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_2.slot_uop_prs1 = 7'b1111111;
    UUT.wrapper.uut.core.int_issue_unit.slots_2.slot_uop_prs2 = 7'b1111111;
    UUT.wrapper.uut.core.int_issue_unit.slots_2.slot_uop_prs3 = 7'b1111111;
    UUT.wrapper.uut.core.int_issue_unit.slots_2.slot_uop_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_2.slot_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_2.slot_uop_taken = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_2.slot_uop_uopc = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_2.slot_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_2.state = 2'b10;
    UUT.wrapper.uut.core.int_issue_unit.slots_3.p1 = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_3.p1_poisoned = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_3.p2 = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_3.p2_poisoned = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_3.p3 = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_3.ppred = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_3.slot_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_3.slot_uop_br_tag = 4'b1111;
    UUT.wrapper.uut.core.int_issue_unit.slots_3.slot_uop_bypassable = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_3.slot_uop_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_3.slot_uop_edge_inst = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_3.slot_uop_ftq_idx = 3'b111;
    UUT.wrapper.uut.core.int_issue_unit.slots_3.slot_uop_fu_code = 10'b0000000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_3.slot_uop_imm_packed = 20'b11111111111111111111;
    UUT.wrapper.uut.core.int_issue_unit.slots_3.slot_uop_is_amo = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_3.slot_uop_is_br = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_3.slot_uop_is_jal = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_3.slot_uop_is_jalr = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_3.slot_uop_is_rvc = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_3.slot_uop_is_sfb = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_3.slot_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_3.slot_uop_ldst_val = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_3.slot_uop_lrs1_rtype = 2'b11;
    UUT.wrapper.uut.core.int_issue_unit.slots_3.slot_uop_lrs2_rtype = 2'b11;
    UUT.wrapper.uut.core.int_issue_unit.slots_3.slot_uop_mem_cmd = 5'b11111;
    UUT.wrapper.uut.core.int_issue_unit.slots_3.slot_uop_pc_lob = 6'b111111;
    UUT.wrapper.uut.core.int_issue_unit.slots_3.slot_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_3.slot_uop_prs1 = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_3.slot_uop_prs2 = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_3.slot_uop_prs3 = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_3.slot_uop_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_3.slot_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_3.slot_uop_taken = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_3.slot_uop_uopc = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_3.slot_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_3.state = 2'b10;
    UUT.wrapper.uut.core.int_issue_unit.slots_4.p1 = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_4.p1_poisoned = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_4.p2 = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_4.p2_poisoned = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_4.p3 = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_4.ppred = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_4.slot_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_4.slot_uop_br_tag = 4'b1111;
    UUT.wrapper.uut.core.int_issue_unit.slots_4.slot_uop_bypassable = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_4.slot_uop_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_4.slot_uop_edge_inst = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_4.slot_uop_ftq_idx = 3'b111;
    UUT.wrapper.uut.core.int_issue_unit.slots_4.slot_uop_fu_code = 10'b0000000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_4.slot_uop_imm_packed = 20'b11111111111111111111;
    UUT.wrapper.uut.core.int_issue_unit.slots_4.slot_uop_is_amo = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_4.slot_uop_is_br = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_4.slot_uop_is_jal = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_4.slot_uop_is_jalr = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_4.slot_uop_is_rvc = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_4.slot_uop_is_sfb = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_4.slot_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_4.slot_uop_ldst_val = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_4.slot_uop_lrs1_rtype = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_4.slot_uop_lrs2_rtype = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_4.slot_uop_mem_cmd = 5'b11111;
    UUT.wrapper.uut.core.int_issue_unit.slots_4.slot_uop_pc_lob = 6'b111111;
    UUT.wrapper.uut.core.int_issue_unit.slots_4.slot_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_4.slot_uop_prs1 = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_4.slot_uop_prs2 = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_4.slot_uop_prs3 = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_4.slot_uop_rob_idx = 6'b111111;
    UUT.wrapper.uut.core.int_issue_unit.slots_4.slot_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_4.slot_uop_taken = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_4.slot_uop_uopc = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_4.slot_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_4.state = 2'b10;
    UUT.wrapper.uut.core.int_issue_unit.slots_5.p1 = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_5.p1_poisoned = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_5.p2 = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_5.p2_poisoned = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_5.p3 = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_5.ppred = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_5.slot_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_5.slot_uop_br_tag = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_5.slot_uop_bypassable = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_5.slot_uop_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_5.slot_uop_edge_inst = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_5.slot_uop_ftq_idx = 3'b000;
    UUT.wrapper.uut.core.int_issue_unit.slots_5.slot_uop_fu_code = 10'b0000000001;
    UUT.wrapper.uut.core.int_issue_unit.slots_5.slot_uop_imm_packed = 20'b00000000000000000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_5.slot_uop_is_amo = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_5.slot_uop_is_br = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_5.slot_uop_is_jal = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_5.slot_uop_is_jalr = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_5.slot_uop_is_rvc = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_5.slot_uop_is_sfb = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_5.slot_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_5.slot_uop_ldst_val = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_5.slot_uop_lrs1_rtype = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_5.slot_uop_lrs2_rtype = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_5.slot_uop_mem_cmd = 5'b00000;
    UUT.wrapper.uut.core.int_issue_unit.slots_5.slot_uop_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_5.slot_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_5.slot_uop_prs1 = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_5.slot_uop_prs2 = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_5.slot_uop_prs3 = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_5.slot_uop_rob_idx = 6'b111111;
    UUT.wrapper.uut.core.int_issue_unit.slots_5.slot_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_5.slot_uop_taken = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_5.slot_uop_uopc = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_5.slot_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_5.state = 2'b11;
    UUT.wrapper.uut.core.int_issue_unit.slots_6.p1 = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_6.p1_poisoned = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_6.p2 = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_6.p2_poisoned = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_6.p3 = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_6.ppred = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_6.slot_uop_br_mask = 12'b111100010000;
    UUT.wrapper.uut.core.int_issue_unit.slots_6.slot_uop_br_tag = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_6.slot_uop_bypassable = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_6.slot_uop_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_6.slot_uop_edge_inst = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_6.slot_uop_ftq_idx = 3'b000;
    UUT.wrapper.uut.core.int_issue_unit.slots_6.slot_uop_fu_code = 10'b0000001011;
    UUT.wrapper.uut.core.int_issue_unit.slots_6.slot_uop_imm_packed = 20'b00000000000000000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_6.slot_uop_is_amo = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_6.slot_uop_is_br = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_6.slot_uop_is_jal = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_6.slot_uop_is_jalr = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_6.slot_uop_is_rvc = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_6.slot_uop_is_sfb = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_6.slot_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_6.slot_uop_ldst_val = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_6.slot_uop_lrs1_rtype = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_6.slot_uop_lrs2_rtype = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_6.slot_uop_mem_cmd = 5'b00000;
    UUT.wrapper.uut.core.int_issue_unit.slots_6.slot_uop_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_6.slot_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_6.slot_uop_prs1 = 7'b0000010;
    UUT.wrapper.uut.core.int_issue_unit.slots_6.slot_uop_prs2 = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_6.slot_uop_prs3 = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_6.slot_uop_rob_idx = 6'b111111;
    UUT.wrapper.uut.core.int_issue_unit.slots_6.slot_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_6.slot_uop_taken = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_6.slot_uop_uopc = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_6.slot_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_6.state = 2'b01;
    UUT.wrapper.uut.core.int_issue_unit.slots_7.p1 = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_7.p1_poisoned = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_7.p2 = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_7.p2_poisoned = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_7.p3 = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_7.ppred = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_7.slot_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_7.slot_uop_br_tag = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_7.slot_uop_bypassable = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_7.slot_uop_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_7.slot_uop_edge_inst = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_7.slot_uop_ftq_idx = 3'b000;
    UUT.wrapper.uut.core.int_issue_unit.slots_7.slot_uop_fu_code = 10'b0000111011;
    UUT.wrapper.uut.core.int_issue_unit.slots_7.slot_uop_imm_packed = 20'b00000000000000000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_7.slot_uop_is_amo = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_7.slot_uop_is_br = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_7.slot_uop_is_jal = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_7.slot_uop_is_jalr = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_7.slot_uop_is_rvc = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_7.slot_uop_is_sfb = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_7.slot_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_7.slot_uop_ldst_val = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_7.slot_uop_lrs1_rtype = 2'b01;
    UUT.wrapper.uut.core.int_issue_unit.slots_7.slot_uop_lrs2_rtype = 2'b01;
    UUT.wrapper.uut.core.int_issue_unit.slots_7.slot_uop_mem_cmd = 5'b00000;
    UUT.wrapper.uut.core.int_issue_unit.slots_7.slot_uop_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_7.slot_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_7.slot_uop_prs1 = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_7.slot_uop_prs2 = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_7.slot_uop_prs3 = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_7.slot_uop_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_7.slot_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_7.slot_uop_taken = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_7.slot_uop_uopc = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_7.slot_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_7.state = 2'b01;
    UUT.wrapper.uut.core.int_issue_unit.slots_8.p1 = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_8.p1_poisoned = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_8.p2 = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_8.p2_poisoned = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_8.p3 = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_8.ppred = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_8.slot_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_8.slot_uop_br_tag = 4'b0001;
    UUT.wrapper.uut.core.int_issue_unit.slots_8.slot_uop_bypassable = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_8.slot_uop_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_8.slot_uop_edge_inst = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_8.slot_uop_ftq_idx = 3'b000;
    UUT.wrapper.uut.core.int_issue_unit.slots_8.slot_uop_fu_code = 10'b0000100001;
    UUT.wrapper.uut.core.int_issue_unit.slots_8.slot_uop_imm_packed = 20'b00000000000000000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_8.slot_uop_is_amo = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_8.slot_uop_is_br = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_8.slot_uop_is_jal = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_8.slot_uop_is_jalr = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_8.slot_uop_is_rvc = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_8.slot_uop_is_sfb = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_8.slot_uop_ldq_idx = 4'b1111;
    UUT.wrapper.uut.core.int_issue_unit.slots_8.slot_uop_ldst_val = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_8.slot_uop_lrs1_rtype = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_8.slot_uop_lrs2_rtype = 2'b10;
    UUT.wrapper.uut.core.int_issue_unit.slots_8.slot_uop_mem_cmd = 5'b00000;
    UUT.wrapper.uut.core.int_issue_unit.slots_8.slot_uop_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_8.slot_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_8.slot_uop_prs1 = 7'b0001010;
    UUT.wrapper.uut.core.int_issue_unit.slots_8.slot_uop_prs2 = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_8.slot_uop_prs3 = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_8.slot_uop_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_8.slot_uop_stq_idx = 4'b1111;
    UUT.wrapper.uut.core.int_issue_unit.slots_8.slot_uop_taken = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_8.slot_uop_uopc = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_8.slot_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_8.state = 2'b01;
    UUT.wrapper.uut.core.int_issue_unit.slots_9.p1 = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_9.p1_poisoned = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_9.p2 = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_9.p2_poisoned = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_9.p3 = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_9.ppred = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_9.slot_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_9.slot_uop_br_tag = 4'b0000;
    UUT.wrapper.uut.core.int_issue_unit.slots_9.slot_uop_bypassable = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_9.slot_uop_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit.slots_9.slot_uop_edge_inst = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_9.slot_uop_ftq_idx = 3'b000;
    UUT.wrapper.uut.core.int_issue_unit.slots_9.slot_uop_fu_code = 10'b0000111011;
    UUT.wrapper.uut.core.int_issue_unit.slots_9.slot_uop_imm_packed = 20'b00000000000000000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_9.slot_uop_is_amo = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_9.slot_uop_is_br = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_9.slot_uop_is_jal = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_9.slot_uop_is_jalr = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_9.slot_uop_is_rvc = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_9.slot_uop_is_sfb = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_9.slot_uop_ldq_idx = 4'b1111;
    UUT.wrapper.uut.core.int_issue_unit.slots_9.slot_uop_ldst_val = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_9.slot_uop_lrs1_rtype = 2'b01;
    UUT.wrapper.uut.core.int_issue_unit.slots_9.slot_uop_lrs2_rtype = 2'b01;
    UUT.wrapper.uut.core.int_issue_unit.slots_9.slot_uop_mem_cmd = 5'b00000;
    UUT.wrapper.uut.core.int_issue_unit.slots_9.slot_uop_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_9.slot_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_9.slot_uop_prs1 = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_9.slot_uop_prs2 = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_9.slot_uop_prs3 = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_9.slot_uop_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_9.slot_uop_stq_idx = 4'b1111;
    UUT.wrapper.uut.core.int_issue_unit.slots_9.slot_uop_taken = 1'b1;
    UUT.wrapper.uut.core.int_issue_unit.slots_9.slot_uop_uopc = 7'b0000000;
    UUT.wrapper.uut.core.int_issue_unit.slots_9.slot_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.core.int_issue_unit.slots_9.state = 2'b00;
    UUT.wrapper.uut.core.int_issue_unit_io_flush_pipeline_REG = 1'b1;
    UUT.wrapper.uut.core.int_regfile_state_0 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.int_regfile_state_1 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.int_regfile_state_10 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.int_regfile_state_11 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.int_regfile_state_12 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.int_regfile_state_13 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.int_regfile_state_14 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.int_regfile_state_15 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.int_regfile_state_16 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.int_regfile_state_17 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.int_regfile_state_18 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.int_regfile_state_19 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.int_regfile_state_2 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.int_regfile_state_20 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.int_regfile_state_21 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.int_regfile_state_22 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.int_regfile_state_23 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.int_regfile_state_24 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.int_regfile_state_25 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.int_regfile_state_26 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.int_regfile_state_27 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.int_regfile_state_28 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.int_regfile_state_29 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.int_regfile_state_3 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.int_regfile_state_30 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.int_regfile_state_31 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.int_regfile_state_4 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.int_regfile_state_5 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.int_regfile_state_6 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.int_regfile_state_7 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.int_regfile_state_8 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.int_regfile_state_9 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.io_ifu_commit_bits_REG = 3'b011;
    UUT.wrapper.uut.core.io_ifu_redirect_ftq_idx_REG = 3'b000;
    UUT.wrapper.uut.core.io_ifu_redirect_pc_REG = 40'b1000000000010000000000000000000000000000;
    UUT.wrapper.uut.core.io_ifu_redirect_pc_REG_1 = 40'b0011111100000000000000000000000000000110;
    UUT.wrapper.uut.core.io_ifu_sfence_REG_bits_addr = 39'b100000100000000000000001111111110000000;
    UUT.wrapper.uut.core.io_ifu_sfence_REG_bits_rs1 = 1'b0;
    UUT.wrapper.uut.core.io_ifu_sfence_REG_bits_rs2 = 1'b0;
    UUT.wrapper.uut.core.io_ifu_sfence_REG_valid = 1'b0;
    UUT.wrapper.uut.core.io_lsu_exception_REG = 1'b0;
    UUT.wrapper.uut.core.iregfile.read_addrs_0 = 7'b0000000;
    UUT.wrapper.uut.core.iregfile.read_addrs_1 = 7'b0000000;
    UUT.wrapper.uut.core.iregfile.read_addrs_2 = 7'b0000000;
    UUT.wrapper.uut.core.iregfile.read_addrs_3 = 7'b0000000;
    UUT.wrapper.uut.core.iregfile.read_addrs_4 = 7'b0000000;
    UUT.wrapper.uut.core.iregfile.read_addrs_5 = 7'b0000000;
    UUT.wrapper.uut.core.iregfile.regfile_0 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_1 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_10 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_11 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_12 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_13 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_14 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_15 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_16 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_17 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_18 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_19 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_2 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_20 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_21 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_22 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_23 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_24 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_25 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_26 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_27 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_28 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_29 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_3 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_30 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_31 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_32 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_33 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_34 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_35 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_36 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_37 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_38 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_39 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_4 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_40 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_41 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_42 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_43 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_44 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_45 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_46 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_47 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_48 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_49 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_5 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_50 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_51 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_52 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_53 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_54 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_55 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_56 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_57 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_58 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_59 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_6 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_60 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_61 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_62 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_63 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_64 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_65 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_66 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_67 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_68 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_69 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_7 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_70 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_71 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_72 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_75 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_78 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_8 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregfile.regfile_9 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregister_read.exe_reg_rs1_data_0 = 64'b0000000000000000000000000001100111111111111111111111000000001100;
    UUT.wrapper.uut.core.iregister_read.exe_reg_rs1_data_1 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregister_read.exe_reg_rs1_data_2 = 64'b1011001110110011001100110011000000000000000000000000000000000001;
    UUT.wrapper.uut.core.iregister_read.exe_reg_rs2_data_0 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregister_read.exe_reg_rs2_data_1 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.iregister_read.exe_reg_rs2_data_2 = 64'b1000000000000000000000000000000000000000000000000000000000000110;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_0_br_mask = 12'b111111111111;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_0_ctrl_is_load = 1'b1;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_0_ctrl_is_sta = 1'b0;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_0_ctrl_is_std = 1'b0;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_0_fp_val = 1'b0;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_0_fu_code = 10'b0000000111;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_0_imm_packed = 20'b10011100110011111111;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_0_is_amo = 1'b0;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_0_ldq_idx = 4'b1100;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_0_mem_cmd = 5'b11000;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_0_mem_signed = 1'b0;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_0_mem_size = 2'b11;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_0_pdst = 7'b0000000;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_0_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_0_stq_idx = 4'b1111;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_0_uopc = 7'b0000000;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_0_uses_ldq = 1'b0;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_0_uses_stq = 1'b0;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_1_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_1_br_tag = 4'b0000;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_1_bypassable = 1'b0;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_1_ctrl_br_type = 4'b0000;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_1_ctrl_fcn_dw = 1'b1;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_1_ctrl_imm_sel = 3'b000;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_1_ctrl_op1_sel = 2'b00;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_1_ctrl_op2_sel = 3'b000;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_1_ctrl_op_fcn = 5'b00011;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_1_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_1_edge_inst = 1'b0;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_1_ftq_idx = 3'b000;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_1_fu_code = 10'b1111111111;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_1_imm_packed = 20'b00000000000000000000;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_1_is_amo = 1'b0;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_1_is_br = 1'b0;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_1_is_jal = 1'b0;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_1_is_jalr = 1'b0;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_1_is_rvc = 1'b0;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_1_is_sfb = 1'b0;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_1_ldq_idx = 4'b0000;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_1_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_1_pdst = 7'b0000000;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_1_prs1 = 7'b0000000;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_1_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_1_stq_idx = 4'b0000;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_1_taken = 1'b0;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_1_uopc = 7'b0000000;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_1_uses_stq = 1'b0;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_2_br_mask = 12'b111111111111;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_2_br_tag = 4'b0000;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_2_bypassable = 1'b0;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_2_ctrl_br_type = 4'b0000;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_2_ctrl_csr_cmd = 3'b000;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_2_ctrl_fcn_dw = 1'b0;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_2_ctrl_imm_sel = 3'b000;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_2_ctrl_op1_sel = 2'b00;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_2_ctrl_op2_sel = 3'b000;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_2_ctrl_op_fcn = 5'b11000;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_2_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_2_edge_inst = 1'b0;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_2_ftq_idx = 3'b000;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_2_fu_code = 10'b1111111111;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_2_imm_packed = 20'b00000000000000000000;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_2_is_amo = 1'b0;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_2_is_br = 1'b0;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_2_is_jal = 1'b0;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_2_is_jalr = 1'b0;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_2_is_rvc = 1'b0;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_2_is_sfb = 1'b0;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_2_ldq_idx = 4'b0000;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_2_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_2_pdst = 7'b0000000;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_2_prs1 = 7'b0000000;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_2_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_2_stq_idx = 4'b0000;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_2_taken = 1'b0;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_2_uopc = 7'b0000000;
    UUT.wrapper.uut.core.iregister_read.exe_reg_uops_2_uses_stq = 1'b0;
    UUT.wrapper.uut.core.iregister_read.exe_reg_valids_0 = 1'b1;
    UUT.wrapper.uut.core.iregister_read.exe_reg_valids_1 = 1'b1;
    UUT.wrapper.uut.core.iregister_read.exe_reg_valids_2 = 1'b0;
    UUT.wrapper.uut.core.iregister_read.rrd_rs1_data_0_REG = 1'b0;
    UUT.wrapper.uut.core.iregister_read.rrd_rs1_data_1_REG = 1'b0;
    UUT.wrapper.uut.core.iregister_read.rrd_rs1_data_2_REG = 1'b0;
    UUT.wrapper.uut.core.iregister_read.rrd_rs2_data_0_REG = 1'b0;
    UUT.wrapper.uut.core.iregister_read.rrd_rs2_data_1_REG = 1'b0;
    UUT.wrapper.uut.core.iregister_read.rrd_rs2_data_2_REG = 1'b0;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_0_REG_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_0_REG_ctrl_is_load = 1'b0;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_0_REG_ctrl_is_sta = 1'b0;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_0_REG_ctrl_is_std = 1'b0;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_0_REG_fp_val = 1'b0;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_0_REG_fu_code = 10'b0000000000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_0_REG_imm_packed = 20'b00000000000000000000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_0_REG_is_amo = 1'b0;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_0_REG_ldq_idx = 4'b0000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_0_REG_lrs1_rtype = 2'b00;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_0_REG_lrs2_rtype = 2'b00;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_0_REG_mem_cmd = 5'b00000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_0_REG_mem_signed = 1'b0;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_0_REG_mem_size = 2'b00;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_0_REG_pdst = 7'b0000000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_0_REG_prs1 = 7'b0000000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_0_REG_prs2 = 7'b0000000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_0_REG_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_0_REG_stq_idx = 4'b0000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_0_REG_uopc = 7'b0000000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_0_REG_uses_ldq = 1'b0;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_0_REG_uses_stq = 1'b0;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_1_REG_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_1_REG_br_tag = 4'b0000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_1_REG_bypassable = 1'b0;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_1_REG_ctrl_br_type = 4'b0000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_1_REG_ctrl_fcn_dw = 1'b0;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_1_REG_ctrl_imm_sel = 3'b000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_1_REG_ctrl_op1_sel = 2'b00;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_1_REG_ctrl_op2_sel = 3'b000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_1_REG_ctrl_op_fcn = 5'b00000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_1_REG_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_1_REG_edge_inst = 1'b0;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_1_REG_ftq_idx = 3'b000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_1_REG_fu_code = 10'b0000000000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_1_REG_imm_packed = 20'b00000000000000000000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_1_REG_is_amo = 1'b0;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_1_REG_is_br = 1'b0;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_1_REG_is_jal = 1'b0;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_1_REG_is_jalr = 1'b0;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_1_REG_is_rvc = 1'b0;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_1_REG_is_sfb = 1'b0;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_1_REG_ldq_idx = 4'b0000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_1_REG_lrs1_rtype = 2'b00;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_1_REG_lrs2_rtype = 2'b00;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_1_REG_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_1_REG_pdst = 7'b0000000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_1_REG_prs1 = 7'b0000000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_1_REG_prs2 = 7'b0000000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_1_REG_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_1_REG_stq_idx = 4'b0000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_1_REG_taken = 1'b0;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_1_REG_uopc = 7'b0000000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_1_REG_uses_stq = 1'b0;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_2_REG_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_2_REG_br_tag = 4'b0000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_2_REG_bypassable = 1'b0;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_2_REG_ctrl_br_type = 4'b0000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_2_REG_ctrl_csr_cmd = 3'b000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_2_REG_ctrl_fcn_dw = 1'b0;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_2_REG_ctrl_imm_sel = 3'b000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_2_REG_ctrl_op1_sel = 2'b00;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_2_REG_ctrl_op2_sel = 3'b000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_2_REG_ctrl_op_fcn = 5'b00000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_2_REG_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_2_REG_edge_inst = 1'b0;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_2_REG_ftq_idx = 3'b000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_2_REG_fu_code = 10'b0000000000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_2_REG_imm_packed = 20'b00000000000000000000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_2_REG_is_amo = 1'b0;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_2_REG_is_br = 1'b0;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_2_REG_is_jal = 1'b0;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_2_REG_is_jalr = 1'b0;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_2_REG_is_rvc = 1'b0;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_2_REG_is_sfb = 1'b0;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_2_REG_ldq_idx = 4'b0000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_2_REG_lrs1_rtype = 2'b00;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_2_REG_lrs2_rtype = 2'b00;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_2_REG_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_2_REG_pdst = 7'b0000000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_2_REG_prs1 = 7'b0000000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_2_REG_prs2 = 7'b0000000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_2_REG_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_2_REG_stq_idx = 4'b0000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_2_REG_taken = 1'b0;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_2_REG_uopc = 7'b0000000;
    UUT.wrapper.uut.core.iregister_read.rrd_uops_2_REG_uses_stq = 1'b0;
    UUT.wrapper.uut.core.iregister_read.rrd_valids_0_REG = 1'b0;
    UUT.wrapper.uut.core.iregister_read.rrd_valids_1_REG = 1'b0;
    UUT.wrapper.uut.core.iregister_read.rrd_valids_2_REG = 1'b0;
    UUT.wrapper.uut.core.iregister_read_io_kill_REG = 1'b0;
    UUT.wrapper.uut.core.jmp_pc_req_bits_REG = 3'b000;
    UUT.wrapper.uut.core.jmp_pc_req_valid_REG = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.io_dis_uops_0_ready_REG = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.io_dis_uops_1_ready_REG = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_0.p1 = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_0.p1_poisoned = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_0.p2 = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_0.p2_poisoned = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_0.p3 = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_0.ppred = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_0.slot_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_0.slot_uop_fp_val = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_0.slot_uop_fu_code = 10'b1111111011;
    UUT.wrapper.uut.core.mem_issue_unit.slots_0.slot_uop_imm_packed = 20'b00000000000011111111;
    UUT.wrapper.uut.core.mem_issue_unit.slots_0.slot_uop_is_amo = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_0.slot_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_0.slot_uop_lrs1_rtype = 2'b00;
    UUT.wrapper.uut.core.mem_issue_unit.slots_0.slot_uop_lrs2_rtype = 2'b00;
    UUT.wrapper.uut.core.mem_issue_unit.slots_0.slot_uop_mem_cmd = 5'b00000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_0.slot_uop_mem_signed = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_0.slot_uop_mem_size = 2'b00;
    UUT.wrapper.uut.core.mem_issue_unit.slots_0.slot_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_0.slot_uop_prs1 = 7'b0000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_0.slot_uop_prs2 = 7'b0000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_0.slot_uop_prs3 = 7'b0000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_0.slot_uop_rob_idx = 6'b111111;
    UUT.wrapper.uut.core.mem_issue_unit.slots_0.slot_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_0.slot_uop_uopc = 7'b0000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_0.slot_uop_uses_ldq = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_0.slot_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_0.state = 2'b10;
    UUT.wrapper.uut.core.mem_issue_unit.slots_1.p1 = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_1.p1_poisoned = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_1.p2 = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_1.p2_poisoned = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_1.p3 = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_1.ppred = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_1.slot_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_1.slot_uop_fp_val = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_1.slot_uop_fu_code = 10'b1111111011;
    UUT.wrapper.uut.core.mem_issue_unit.slots_1.slot_uop_imm_packed = 20'b00000000000011111111;
    UUT.wrapper.uut.core.mem_issue_unit.slots_1.slot_uop_is_amo = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_1.slot_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_1.slot_uop_lrs1_rtype = 2'b00;
    UUT.wrapper.uut.core.mem_issue_unit.slots_1.slot_uop_lrs2_rtype = 2'b10;
    UUT.wrapper.uut.core.mem_issue_unit.slots_1.slot_uop_mem_cmd = 5'b00000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_1.slot_uop_mem_signed = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_1.slot_uop_mem_size = 2'b00;
    UUT.wrapper.uut.core.mem_issue_unit.slots_1.slot_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_1.slot_uop_prs1 = 7'b0000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_1.slot_uop_prs2 = 7'b0000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_1.slot_uop_prs3 = 7'b1000001;
    UUT.wrapper.uut.core.mem_issue_unit.slots_1.slot_uop_rob_idx = 6'b111111;
    UUT.wrapper.uut.core.mem_issue_unit.slots_1.slot_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_1.slot_uop_uopc = 7'b0000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_1.slot_uop_uses_ldq = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_1.slot_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_1.state = 2'b00;
    UUT.wrapper.uut.core.mem_issue_unit.slots_10.p1 = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_10.p1_poisoned = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_10.p2 = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_10.p2_poisoned = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_10.p3 = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_10.ppred = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_10.slot_uop_br_mask = 12'b001100000001;
    UUT.wrapper.uut.core.mem_issue_unit.slots_10.slot_uop_fp_val = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_10.slot_uop_fu_code = 10'b0000000100;
    UUT.wrapper.uut.core.mem_issue_unit.slots_10.slot_uop_imm_packed = 20'b00000000000000000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_10.slot_uop_is_amo = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_10.slot_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_10.slot_uop_lrs1_rtype = 2'b00;
    UUT.wrapper.uut.core.mem_issue_unit.slots_10.slot_uop_lrs2_rtype = 2'b00;
    UUT.wrapper.uut.core.mem_issue_unit.slots_10.slot_uop_mem_cmd = 5'b00000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_10.slot_uop_mem_signed = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_10.slot_uop_mem_size = 2'b00;
    UUT.wrapper.uut.core.mem_issue_unit.slots_10.slot_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_10.slot_uop_prs1 = 7'b0000010;
    UUT.wrapper.uut.core.mem_issue_unit.slots_10.slot_uop_prs2 = 7'b0000010;
    UUT.wrapper.uut.core.mem_issue_unit.slots_10.slot_uop_prs3 = 7'b0000001;
    UUT.wrapper.uut.core.mem_issue_unit.slots_10.slot_uop_rob_idx = 6'b000011;
    UUT.wrapper.uut.core.mem_issue_unit.slots_10.slot_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_10.slot_uop_uopc = 7'b0000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_10.slot_uop_uses_ldq = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_10.slot_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_10.state = 2'b00;
    UUT.wrapper.uut.core.mem_issue_unit.slots_11.p1 = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_11.p1_poisoned = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_11.p2 = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_11.p2_poisoned = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_11.p3 = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_11.ppred = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_11.slot_uop_br_mask = 12'b000000000010;
    UUT.wrapper.uut.core.mem_issue_unit.slots_11.slot_uop_fp_val = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_11.slot_uop_fu_code = 10'b0000000100;
    UUT.wrapper.uut.core.mem_issue_unit.slots_11.slot_uop_imm_packed = 20'b00110010000000000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_11.slot_uop_is_amo = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_11.slot_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_11.slot_uop_lrs1_rtype = 2'b00;
    UUT.wrapper.uut.core.mem_issue_unit.slots_11.slot_uop_lrs2_rtype = 2'b00;
    UUT.wrapper.uut.core.mem_issue_unit.slots_11.slot_uop_mem_cmd = 5'b00001;
    UUT.wrapper.uut.core.mem_issue_unit.slots_11.slot_uop_mem_signed = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_11.slot_uop_mem_size = 2'b01;
    UUT.wrapper.uut.core.mem_issue_unit.slots_11.slot_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_11.slot_uop_prs1 = 7'b0000001;
    UUT.wrapper.uut.core.mem_issue_unit.slots_11.slot_uop_prs2 = 7'b1000001;
    UUT.wrapper.uut.core.mem_issue_unit.slots_11.slot_uop_prs3 = 7'b0000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_11.slot_uop_rob_idx = 6'b000011;
    UUT.wrapper.uut.core.mem_issue_unit.slots_11.slot_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_11.slot_uop_uopc = 7'b0000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_11.slot_uop_uses_ldq = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_11.slot_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_11.state = 2'b00;
    UUT.wrapper.uut.core.mem_issue_unit.slots_2.p1 = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_2.p1_poisoned = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_2.p2 = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_2.p2_poisoned = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_2.p3 = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_2.ppred = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_2.slot_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_2.slot_uop_fp_val = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_2.slot_uop_fu_code = 10'b1111111111;
    UUT.wrapper.uut.core.mem_issue_unit.slots_2.slot_uop_imm_packed = 20'b00000000000011111111;
    UUT.wrapper.uut.core.mem_issue_unit.slots_2.slot_uop_is_amo = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_2.slot_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_2.slot_uop_lrs1_rtype = 2'b00;
    UUT.wrapper.uut.core.mem_issue_unit.slots_2.slot_uop_lrs2_rtype = 2'b10;
    UUT.wrapper.uut.core.mem_issue_unit.slots_2.slot_uop_mem_cmd = 5'b10100;
    UUT.wrapper.uut.core.mem_issue_unit.slots_2.slot_uop_mem_signed = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_2.slot_uop_mem_size = 2'b00;
    UUT.wrapper.uut.core.mem_issue_unit.slots_2.slot_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_2.slot_uop_prs1 = 7'b0000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_2.slot_uop_prs2 = 7'b0000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_2.slot_uop_prs3 = 7'b0000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_2.slot_uop_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_2.slot_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_2.slot_uop_uopc = 7'b0000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_2.slot_uop_uses_ldq = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_2.slot_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_2.state = 2'b00;
    UUT.wrapper.uut.core.mem_issue_unit.slots_3.p1 = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_3.p1_poisoned = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_3.p2 = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_3.p2_poisoned = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_3.p3 = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_3.ppred = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_3.slot_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_3.slot_uop_fp_val = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_3.slot_uop_fu_code = 10'b1111111111;
    UUT.wrapper.uut.core.mem_issue_unit.slots_3.slot_uop_imm_packed = 20'b00000000000011111111;
    UUT.wrapper.uut.core.mem_issue_unit.slots_3.slot_uop_is_amo = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_3.slot_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_3.slot_uop_lrs1_rtype = 2'b00;
    UUT.wrapper.uut.core.mem_issue_unit.slots_3.slot_uop_lrs2_rtype = 2'b10;
    UUT.wrapper.uut.core.mem_issue_unit.slots_3.slot_uop_mem_cmd = 5'b00000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_3.slot_uop_mem_signed = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_3.slot_uop_mem_size = 2'b00;
    UUT.wrapper.uut.core.mem_issue_unit.slots_3.slot_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_3.slot_uop_prs1 = 7'b0000001;
    UUT.wrapper.uut.core.mem_issue_unit.slots_3.slot_uop_prs2 = 7'b0000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_3.slot_uop_prs3 = 7'b0000010;
    UUT.wrapper.uut.core.mem_issue_unit.slots_3.slot_uop_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_3.slot_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_3.slot_uop_uopc = 7'b0000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_3.slot_uop_uses_ldq = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_3.slot_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_3.state = 2'b00;
    UUT.wrapper.uut.core.mem_issue_unit.slots_4.p1 = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_4.p1_poisoned = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_4.p2 = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_4.p2_poisoned = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_4.p3 = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_4.ppred = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_4.slot_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_4.slot_uop_fp_val = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_4.slot_uop_fu_code = 10'b0000010110;
    UUT.wrapper.uut.core.mem_issue_unit.slots_4.slot_uop_imm_packed = 20'b00000000000011111111;
    UUT.wrapper.uut.core.mem_issue_unit.slots_4.slot_uop_is_amo = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_4.slot_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_4.slot_uop_lrs1_rtype = 2'b01;
    UUT.wrapper.uut.core.mem_issue_unit.slots_4.slot_uop_lrs2_rtype = 2'b01;
    UUT.wrapper.uut.core.mem_issue_unit.slots_4.slot_uop_mem_cmd = 5'b00001;
    UUT.wrapper.uut.core.mem_issue_unit.slots_4.slot_uop_mem_signed = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_4.slot_uop_mem_size = 2'b00;
    UUT.wrapper.uut.core.mem_issue_unit.slots_4.slot_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_4.slot_uop_prs1 = 7'b0000010;
    UUT.wrapper.uut.core.mem_issue_unit.slots_4.slot_uop_prs2 = 7'b0000010;
    UUT.wrapper.uut.core.mem_issue_unit.slots_4.slot_uop_prs3 = 7'b0000010;
    UUT.wrapper.uut.core.mem_issue_unit.slots_4.slot_uop_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_4.slot_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_4.slot_uop_uopc = 7'b0000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_4.slot_uop_uses_ldq = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_4.slot_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_4.state = 2'b00;
    UUT.wrapper.uut.core.mem_issue_unit.slots_5.p1 = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_5.p1_poisoned = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_5.p2 = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_5.p2_poisoned = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_5.p3 = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_5.ppred = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_5.slot_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_5.slot_uop_fp_val = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_5.slot_uop_fu_code = 10'b0000010110;
    UUT.wrapper.uut.core.mem_issue_unit.slots_5.slot_uop_imm_packed = 20'b00000000000011111111;
    UUT.wrapper.uut.core.mem_issue_unit.slots_5.slot_uop_is_amo = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_5.slot_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_5.slot_uop_lrs1_rtype = 2'b10;
    UUT.wrapper.uut.core.mem_issue_unit.slots_5.slot_uop_lrs2_rtype = 2'b00;
    UUT.wrapper.uut.core.mem_issue_unit.slots_5.slot_uop_mem_cmd = 5'b00001;
    UUT.wrapper.uut.core.mem_issue_unit.slots_5.slot_uop_mem_signed = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_5.slot_uop_mem_size = 2'b00;
    UUT.wrapper.uut.core.mem_issue_unit.slots_5.slot_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_5.slot_uop_prs1 = 7'b0000001;
    UUT.wrapper.uut.core.mem_issue_unit.slots_5.slot_uop_prs2 = 7'b0000111;
    UUT.wrapper.uut.core.mem_issue_unit.slots_5.slot_uop_prs3 = 7'b0000001;
    UUT.wrapper.uut.core.mem_issue_unit.slots_5.slot_uop_rob_idx = 6'b000001;
    UUT.wrapper.uut.core.mem_issue_unit.slots_5.slot_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_5.slot_uop_uopc = 7'b0000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_5.slot_uop_uses_ldq = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_5.slot_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_5.state = 2'b00;
    UUT.wrapper.uut.core.mem_issue_unit.slots_6.p1 = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_6.p1_poisoned = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_6.p2 = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_6.p2_poisoned = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_6.p3 = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_6.ppred = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_6.slot_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_6.slot_uop_fp_val = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_6.slot_uop_fu_code = 10'b0000010110;
    UUT.wrapper.uut.core.mem_issue_unit.slots_6.slot_uop_imm_packed = 20'b00000000000011111111;
    UUT.wrapper.uut.core.mem_issue_unit.slots_6.slot_uop_is_amo = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_6.slot_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_6.slot_uop_lrs1_rtype = 2'b01;
    UUT.wrapper.uut.core.mem_issue_unit.slots_6.slot_uop_lrs2_rtype = 2'b10;
    UUT.wrapper.uut.core.mem_issue_unit.slots_6.slot_uop_mem_cmd = 5'b00001;
    UUT.wrapper.uut.core.mem_issue_unit.slots_6.slot_uop_mem_signed = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_6.slot_uop_mem_size = 2'b00;
    UUT.wrapper.uut.core.mem_issue_unit.slots_6.slot_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_6.slot_uop_prs1 = 7'b0000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_6.slot_uop_prs2 = 7'b0001001;
    UUT.wrapper.uut.core.mem_issue_unit.slots_6.slot_uop_prs3 = 7'b0000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_6.slot_uop_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_6.slot_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_6.slot_uop_uopc = 7'b0000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_6.slot_uop_uses_ldq = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_6.slot_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_6.state = 2'b00;
    UUT.wrapper.uut.core.mem_issue_unit.slots_7.p1 = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_7.p1_poisoned = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_7.p2 = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_7.p2_poisoned = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_7.p3 = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_7.ppred = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_7.slot_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_7.slot_uop_fp_val = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_7.slot_uop_fu_code = 10'b0000000101;
    UUT.wrapper.uut.core.mem_issue_unit.slots_7.slot_uop_imm_packed = 20'b01111101010011111111;
    UUT.wrapper.uut.core.mem_issue_unit.slots_7.slot_uop_is_amo = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_7.slot_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_7.slot_uop_lrs1_rtype = 2'b00;
    UUT.wrapper.uut.core.mem_issue_unit.slots_7.slot_uop_lrs2_rtype = 2'b00;
    UUT.wrapper.uut.core.mem_issue_unit.slots_7.slot_uop_mem_cmd = 5'b00001;
    UUT.wrapper.uut.core.mem_issue_unit.slots_7.slot_uop_mem_signed = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_7.slot_uop_mem_size = 2'b00;
    UUT.wrapper.uut.core.mem_issue_unit.slots_7.slot_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_7.slot_uop_prs1 = 7'b0010000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_7.slot_uop_prs2 = 7'b1000011;
    UUT.wrapper.uut.core.mem_issue_unit.slots_7.slot_uop_prs3 = 7'b0000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_7.slot_uop_rob_idx = 6'b000011;
    UUT.wrapper.uut.core.mem_issue_unit.slots_7.slot_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_7.slot_uop_uopc = 7'b0000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_7.slot_uop_uses_ldq = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_7.slot_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_7.state = 2'b00;
    UUT.wrapper.uut.core.mem_issue_unit.slots_8.p1 = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_8.p1_poisoned = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_8.p2 = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_8.p2_poisoned = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_8.p3 = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_8.ppred = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_8.slot_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_8.slot_uop_fp_val = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_8.slot_uop_fu_code = 10'b0000000101;
    UUT.wrapper.uut.core.mem_issue_unit.slots_8.slot_uop_imm_packed = 20'b00000010000000000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_8.slot_uop_is_amo = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_8.slot_uop_ldq_idx = 4'b0001;
    UUT.wrapper.uut.core.mem_issue_unit.slots_8.slot_uop_lrs1_rtype = 2'b01;
    UUT.wrapper.uut.core.mem_issue_unit.slots_8.slot_uop_lrs2_rtype = 2'b10;
    UUT.wrapper.uut.core.mem_issue_unit.slots_8.slot_uop_mem_cmd = 5'b00000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_8.slot_uop_mem_signed = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_8.slot_uop_mem_size = 2'b10;
    UUT.wrapper.uut.core.mem_issue_unit.slots_8.slot_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_8.slot_uop_prs1 = 7'b1000011;
    UUT.wrapper.uut.core.mem_issue_unit.slots_8.slot_uop_prs2 = 7'b1000001;
    UUT.wrapper.uut.core.mem_issue_unit.slots_8.slot_uop_prs3 = 7'b0000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_8.slot_uop_rob_idx = 6'b000010;
    UUT.wrapper.uut.core.mem_issue_unit.slots_8.slot_uop_stq_idx = 4'b0001;
    UUT.wrapper.uut.core.mem_issue_unit.slots_8.slot_uop_uopc = 7'b0000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_8.slot_uop_uses_ldq = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_8.slot_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_8.state = 2'b00;
    UUT.wrapper.uut.core.mem_issue_unit.slots_9.p1 = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_9.p1_poisoned = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_9.p2 = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_9.p2_poisoned = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_9.p3 = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_9.ppred = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_9.slot_uop_br_mask = 12'b000000000010;
    UUT.wrapper.uut.core.mem_issue_unit.slots_9.slot_uop_fp_val = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_9.slot_uop_fu_code = 10'b0000000100;
    UUT.wrapper.uut.core.mem_issue_unit.slots_9.slot_uop_imm_packed = 20'b00100001100000000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_9.slot_uop_is_amo = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_9.slot_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_9.slot_uop_lrs1_rtype = 2'b00;
    UUT.wrapper.uut.core.mem_issue_unit.slots_9.slot_uop_lrs2_rtype = 2'b10;
    UUT.wrapper.uut.core.mem_issue_unit.slots_9.slot_uop_mem_cmd = 5'b00001;
    UUT.wrapper.uut.core.mem_issue_unit.slots_9.slot_uop_mem_signed = 1'b1;
    UUT.wrapper.uut.core.mem_issue_unit.slots_9.slot_uop_mem_size = 2'b11;
    UUT.wrapper.uut.core.mem_issue_unit.slots_9.slot_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_9.slot_uop_prs1 = 7'b0000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_9.slot_uop_prs2 = 7'b0000101;
    UUT.wrapper.uut.core.mem_issue_unit.slots_9.slot_uop_prs3 = 7'b0000100;
    UUT.wrapper.uut.core.mem_issue_unit.slots_9.slot_uop_rob_idx = 6'b000001;
    UUT.wrapper.uut.core.mem_issue_unit.slots_9.slot_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_9.slot_uop_uopc = 7'b0000000;
    UUT.wrapper.uut.core.mem_issue_unit.slots_9.slot_uop_uses_ldq = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_9.slot_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.core.mem_issue_unit.slots_9.state = 2'b00;
    UUT.wrapper.uut.core.mem_issue_unit_io_flush_pipeline_REG = 1'b1;
    UUT.wrapper.uut.core.pause_mem_REG = 1'b1;
    UUT.wrapper.uut.core.rename_stage.busytable.busy_table = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rename_stage.freelist.br_alloc_lists_0 = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rename_stage.freelist.br_alloc_lists_1 = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rename_stage.freelist.br_alloc_lists_10 = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rename_stage.freelist.br_alloc_lists_11 = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rename_stage.freelist.br_alloc_lists_2 = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rename_stage.freelist.br_alloc_lists_3 = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rename_stage.freelist.br_alloc_lists_4 = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rename_stage.freelist.br_alloc_lists_5 = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rename_stage.freelist.br_alloc_lists_6 = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rename_stage.freelist.br_alloc_lists_7 = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rename_stage.freelist.br_alloc_lists_8 = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rename_stage.freelist.br_alloc_lists_9 = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rename_stage.freelist.free_list = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rename_stage.freelist.r_sel = 7'b1110000;
    UUT.wrapper.uut.core.rename_stage.freelist.r_sel_1 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.freelist.r_valid = 1'b1;
    UUT.wrapper.uut.core.rename_stage.freelist.r_valid_1 = 1'b1;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_0_1 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_0_10 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_0_11 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_0_12 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_0_13 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_0_14 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_0_15 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_0_16 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_0_17 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_0_18 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_0_19 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_0_2 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_0_20 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_0_21 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_0_22 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_0_23 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_0_24 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_0_25 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_0_26 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_0_27 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_0_28 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_0_29 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_0_3 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_0_30 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_0_31 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_0_4 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_0_5 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_0_6 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_0_7 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_0_8 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_0_9 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_10_1 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_10_10 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_10_11 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_10_12 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_10_13 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_10_14 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_10_15 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_10_16 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_10_17 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_10_18 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_10_19 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_10_2 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_10_20 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_10_21 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_10_22 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_10_23 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_10_24 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_10_25 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_10_26 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_10_27 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_10_28 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_10_29 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_10_3 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_10_30 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_10_31 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_10_4 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_10_5 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_10_6 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_10_7 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_10_8 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_10_9 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_11_1 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_11_10 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_11_11 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_11_12 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_11_13 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_11_14 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_11_15 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_11_16 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_11_17 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_11_18 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_11_19 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_11_2 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_11_20 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_11_21 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_11_22 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_11_23 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_11_24 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_11_25 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_11_26 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_11_27 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_11_28 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_11_29 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_11_3 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_11_30 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_11_31 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_11_4 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_11_5 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_11_6 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_11_7 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_11_8 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_11_9 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_1_1 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_1_10 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_1_11 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_1_12 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_1_13 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_1_14 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_1_15 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_1_16 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_1_17 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_1_18 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_1_19 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_1_2 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_1_20 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_1_21 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_1_22 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_1_23 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_1_24 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_1_25 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_1_26 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_1_27 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_1_28 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_1_29 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_1_3 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_1_30 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_1_31 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_1_4 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_1_5 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_1_6 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_1_7 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_1_8 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_1_9 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_2_1 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_2_10 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_2_11 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_2_12 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_2_13 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_2_14 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_2_15 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_2_16 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_2_17 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_2_18 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_2_19 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_2_2 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_2_20 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_2_21 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_2_22 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_2_23 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_2_24 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_2_25 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_2_26 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_2_27 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_2_28 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_2_29 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_2_3 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_2_30 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_2_31 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_2_4 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_2_5 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_2_6 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_2_7 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_2_8 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_2_9 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_3_1 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_3_10 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_3_11 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_3_12 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_3_13 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_3_14 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_3_15 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_3_16 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_3_17 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_3_18 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_3_19 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_3_2 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_3_20 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_3_21 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_3_22 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_3_23 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_3_24 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_3_25 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_3_26 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_3_27 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_3_28 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_3_29 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_3_3 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_3_30 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_3_31 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_3_4 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_3_5 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_3_6 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_3_7 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_3_8 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_3_9 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_4_1 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_4_10 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_4_11 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_4_12 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_4_13 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_4_14 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_4_15 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_4_16 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_4_17 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_4_18 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_4_19 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_4_2 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_4_20 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_4_21 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_4_22 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_4_23 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_4_24 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_4_25 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_4_26 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_4_27 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_4_28 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_4_29 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_4_3 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_4_30 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_4_31 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_4_4 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_4_5 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_4_6 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_4_7 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_4_8 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_4_9 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_5_1 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_5_10 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_5_11 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_5_12 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_5_13 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_5_14 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_5_15 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_5_16 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_5_17 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_5_18 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_5_19 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_5_2 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_5_20 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_5_21 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_5_22 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_5_23 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_5_24 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_5_25 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_5_26 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_5_27 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_5_28 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_5_29 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_5_3 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_5_30 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_5_31 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_5_4 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_5_5 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_5_6 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_5_7 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_5_8 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_5_9 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_6_1 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_6_10 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_6_11 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_6_12 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_6_13 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_6_14 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_6_15 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_6_16 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_6_17 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_6_18 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_6_19 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_6_2 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_6_20 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_6_21 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_6_22 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_6_23 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_6_24 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_6_25 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_6_26 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_6_27 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_6_28 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_6_29 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_6_3 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_6_30 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_6_31 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_6_4 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_6_5 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_6_6 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_6_7 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_6_8 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_6_9 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_7_1 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_7_10 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_7_11 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_7_12 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_7_13 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_7_14 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_7_15 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_7_16 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_7_17 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_7_18 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_7_19 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_7_2 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_7_20 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_7_21 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_7_22 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_7_23 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_7_24 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_7_25 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_7_26 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_7_27 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_7_28 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_7_29 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_7_3 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_7_30 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_7_31 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_7_4 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_7_5 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_7_6 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_7_7 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_7_8 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_7_9 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_8_1 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_8_10 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_8_11 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_8_12 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_8_13 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_8_14 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_8_15 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_8_16 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_8_17 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_8_18 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_8_19 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_8_2 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_8_20 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_8_21 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_8_22 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_8_23 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_8_24 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_8_25 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_8_26 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_8_27 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_8_28 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_8_29 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_8_3 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_8_30 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_8_31 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_8_4 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_8_5 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_8_6 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_8_7 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_8_8 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_8_9 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_9_1 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_9_10 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_9_11 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_9_12 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_9_13 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_9_14 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_9_15 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_9_16 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_9_17 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_9_18 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_9_19 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_9_2 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_9_20 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_9_21 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_9_22 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_9_23 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_9_24 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_9_25 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_9_26 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_9_27 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_9_28 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_9_29 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_9_3 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_9_30 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_9_31 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_9_4 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_9_5 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_9_6 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_9_7 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_9_8 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.br_snapshots_9_9 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.map_table_1 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.map_table_10 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.map_table_11 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.map_table_12 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.map_table_13 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.map_table_14 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.map_table_15 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.map_table_16 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.map_table_17 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.map_table_18 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.map_table_19 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.map_table_2 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.map_table_20 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.map_table_21 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.map_table_22 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.map_table_23 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.map_table_24 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.map_table_25 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.map_table_26 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.map_table_27 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.map_table_28 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.map_table_29 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.map_table_3 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.map_table_30 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.map_table_31 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.map_table_4 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.map_table_5 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.map_table_6 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.map_table_7 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.map_table_8 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.maptable.map_table_9 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.r_uop_1_br_mask = 12'b000000000001;
    UUT.wrapper.uut.core.rename_stage.r_uop_1_br_tag = 4'b0000;
    UUT.wrapper.uut.core.rename_stage.r_uop_1_bypassable = 1'b0;
    UUT.wrapper.uut.core.rename_stage.r_uop_1_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rename_stage.r_uop_1_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rename_stage.r_uop_1_dst_rtype = 2'b11;
    UUT.wrapper.uut.core.rename_stage.r_uop_1_edge_inst = 1'b0;
    UUT.wrapper.uut.core.rename_stage.r_uop_1_exc_cause = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rename_stage.r_uop_1_exception = 1'b0;
    UUT.wrapper.uut.core.rename_stage.r_uop_1_flush_on_commit = 1'b0;
    UUT.wrapper.uut.core.rename_stage.r_uop_1_fp_val = 1'b0;
    UUT.wrapper.uut.core.rename_stage.r_uop_1_ftq_idx = 3'b000;
    UUT.wrapper.uut.core.rename_stage.r_uop_1_fu_code = 10'b0000000101;
    UUT.wrapper.uut.core.rename_stage.r_uop_1_imm_packed = 20'b00000000000000000000;
    UUT.wrapper.uut.core.rename_stage.r_uop_1_iq_type = 3'b101;
    UUT.wrapper.uut.core.rename_stage.r_uop_1_is_amo = 1'b0;
    UUT.wrapper.uut.core.rename_stage.r_uop_1_is_br = 1'b1;
    UUT.wrapper.uut.core.rename_stage.r_uop_1_is_fence = 1'b0;
    UUT.wrapper.uut.core.rename_stage.r_uop_1_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rename_stage.r_uop_1_is_jal = 1'b1;
    UUT.wrapper.uut.core.rename_stage.r_uop_1_is_jalr = 1'b1;
    UUT.wrapper.uut.core.rename_stage.r_uop_1_is_rvc = 1'b1;
    UUT.wrapper.uut.core.rename_stage.r_uop_1_is_sfb = 1'b1;
    UUT.wrapper.uut.core.rename_stage.r_uop_1_is_sys_pc2epc = 1'b0;
    UUT.wrapper.uut.core.rename_stage.r_uop_1_is_unique = 1'b0;
    UUT.wrapper.uut.core.rename_stage.r_uop_1_ldst = 5'b00001;
    UUT.wrapper.uut.core.rename_stage.r_uop_1_ldst_val = 1'b1;
    UUT.wrapper.uut.core.rename_stage.r_uop_1_lrs1 = 5'b00010;
    UUT.wrapper.uut.core.rename_stage.r_uop_1_lrs1_rtype = 2'b00;
    UUT.wrapper.uut.core.rename_stage.r_uop_1_lrs2 = 5'b10000;
    UUT.wrapper.uut.core.rename_stage.r_uop_1_lrs2_rtype = 2'b01;
    UUT.wrapper.uut.core.rename_stage.r_uop_1_mem_cmd = 5'b00001;
    UUT.wrapper.uut.core.rename_stage.r_uop_1_mem_signed = 1'b1;
    UUT.wrapper.uut.core.rename_stage.r_uop_1_mem_size = 2'b01;
    UUT.wrapper.uut.core.rename_stage.r_uop_1_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.rename_stage.r_uop_1_prs1 = 7'b0000011;
    UUT.wrapper.uut.core.rename_stage.r_uop_1_prs2 = 7'b0000001;
    UUT.wrapper.uut.core.rename_stage.r_uop_1_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.r_uop_1_taken = 1'b1;
    UUT.wrapper.uut.core.rename_stage.r_uop_1_uopc = 7'b0100010;
    UUT.wrapper.uut.core.rename_stage.r_uop_1_uses_ldq = 1'b0;
    UUT.wrapper.uut.core.rename_stage.r_uop_1_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rename_stage.r_uop_br_mask = 12'b010111111110;
    UUT.wrapper.uut.core.rename_stage.r_uop_br_tag = 4'b0000;
    UUT.wrapper.uut.core.rename_stage.r_uop_bypassable = 1'b0;
    UUT.wrapper.uut.core.rename_stage.r_uop_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rename_stage.r_uop_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rename_stage.r_uop_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rename_stage.r_uop_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rename_stage.r_uop_exc_cause = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rename_stage.r_uop_exception = 1'b0;
    UUT.wrapper.uut.core.rename_stage.r_uop_flush_on_commit = 1'b0;
    UUT.wrapper.uut.core.rename_stage.r_uop_fp_val = 1'b0;
    UUT.wrapper.uut.core.rename_stage.r_uop_ftq_idx = 3'b000;
    UUT.wrapper.uut.core.rename_stage.r_uop_fu_code = 10'b0000000100;
    UUT.wrapper.uut.core.rename_stage.r_uop_imm_packed = 20'b11111111111100000000;
    UUT.wrapper.uut.core.rename_stage.r_uop_iq_type = 3'b101;
    UUT.wrapper.uut.core.rename_stage.r_uop_is_amo = 1'b0;
    UUT.wrapper.uut.core.rename_stage.r_uop_is_br = 1'b1;
    UUT.wrapper.uut.core.rename_stage.r_uop_is_fence = 1'b0;
    UUT.wrapper.uut.core.rename_stage.r_uop_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rename_stage.r_uop_is_jal = 1'b1;
    UUT.wrapper.uut.core.rename_stage.r_uop_is_jalr = 1'b1;
    UUT.wrapper.uut.core.rename_stage.r_uop_is_rvc = 1'b1;
    UUT.wrapper.uut.core.rename_stage.r_uop_is_sfb = 1'b1;
    UUT.wrapper.uut.core.rename_stage.r_uop_is_sys_pc2epc = 1'b0;
    UUT.wrapper.uut.core.rename_stage.r_uop_is_unique = 1'b0;
    UUT.wrapper.uut.core.rename_stage.r_uop_ldst = 5'b00000;
    UUT.wrapper.uut.core.rename_stage.r_uop_ldst_val = 1'b1;
    UUT.wrapper.uut.core.rename_stage.r_uop_lrs1 = 5'b11101;
    UUT.wrapper.uut.core.rename_stage.r_uop_lrs1_rtype = 2'b11;
    UUT.wrapper.uut.core.rename_stage.r_uop_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rename_stage.r_uop_lrs2_rtype = 2'b00;
    UUT.wrapper.uut.core.rename_stage.r_uop_mem_cmd = 5'b00000;
    UUT.wrapper.uut.core.rename_stage.r_uop_mem_signed = 1'b0;
    UUT.wrapper.uut.core.rename_stage.r_uop_mem_size = 2'b10;
    UUT.wrapper.uut.core.rename_stage.r_uop_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.rename_stage.r_uop_prs1 = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.r_uop_prs2 = 7'b1111111;
    UUT.wrapper.uut.core.rename_stage.r_uop_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rename_stage.r_uop_taken = 1'b1;
    UUT.wrapper.uut.core.rename_stage.r_uop_uopc = 7'b0100010;
    UUT.wrapper.uut.core.rename_stage.r_uop_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rename_stage.r_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.core.rename_stage.r_valid = 1'b1;
    UUT.wrapper.uut.core.rename_stage.r_valid_1 = 1'b1;
    UUT.wrapper.uut.core.rob.REG = 1'b0;
    UUT.wrapper.uut.core.rob.REG_1 = 1'b0;
    UUT.wrapper.uut.core.rob.REG_2 = 1'b0;
    UUT.wrapper.uut.core.rob.block_commit_REG = 1'b0;
    UUT.wrapper.uut.core.rob.block_commit_REG_1 = 1'b0;
    UUT.wrapper.uut.core.rob.block_commit_REG_2 = 1'b0;
    UUT.wrapper.uut.core.rob.io_com_load_is_at_rob_head_REG = 1'b0;
    UUT.wrapper.uut.core.rob.maybe_full = 1'b0;
    UUT.wrapper.uut.core.rob.r_partial_row = 1'b0;
    UUT.wrapper.uut.core.rob.r_xcpt_badvaddr = 40'b1111111111111111111111111111111111111111;
    UUT.wrapper.uut.core.rob.r_xcpt_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.r_xcpt_uop_exc_cause = 64'b0000000000000000000000000000000000000000000000000000000000010001;
    UUT.wrapper.uut.core.rob.r_xcpt_uop_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.r_xcpt_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_bsy_1_0 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_bsy_1_1 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_bsy_1_10 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_bsy_1_11 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_bsy_1_12 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_bsy_1_13 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_bsy_1_14 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_bsy_1_15 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_bsy_1_16 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_bsy_1_17 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_bsy_1_18 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_bsy_1_19 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_bsy_1_2 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_bsy_1_20 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_bsy_1_21 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_bsy_1_22 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_bsy_1_23 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_bsy_1_24 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_bsy_1_25 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_bsy_1_26 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_bsy_1_27 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_bsy_1_28 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_bsy_1_29 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_bsy_1_3 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_bsy_1_30 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_bsy_1_31 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_bsy_1_4 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_bsy_1_5 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_bsy_1_6 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_bsy_1_7 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_bsy_1_8 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_bsy_1_9 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_bsy__0 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_bsy__1 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_bsy__10 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_bsy__11 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_bsy__12 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_bsy__13 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_bsy__14 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_bsy__15 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_bsy__16 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_bsy__17 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_bsy__18 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_bsy__19 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_bsy__2 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_bsy__20 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_bsy__21 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_bsy__22 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_bsy__23 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_bsy__24 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_bsy__25 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_bsy__26 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_bsy__27 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_bsy__28 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_bsy__29 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_bsy__3 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_bsy__30 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_bsy__31 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_bsy__4 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_bsy__5 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_bsy__6 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_bsy__7 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_bsy__8 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_bsy__9 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_exception_1_0 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_exception_1_1 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_exception_1_10 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_exception_1_11 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_exception_1_12 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_exception_1_13 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_exception_1_14 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_exception_1_15 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_exception_1_16 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_exception_1_17 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_exception_1_18 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_exception_1_19 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_exception_1_2 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_exception_1_20 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_exception_1_21 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_exception_1_22 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_exception_1_23 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_exception_1_24 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_exception_1_25 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_exception_1_26 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_exception_1_27 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_exception_1_28 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_exception_1_29 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_exception_1_3 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_exception_1_30 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_exception_1_31 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_exception_1_4 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_exception_1_5 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_exception_1_6 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_exception_1_7 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_exception_1_8 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_exception_1_9 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_exception__0 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_exception__1 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_exception__10 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_exception__11 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_exception__12 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_exception__13 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_exception__14 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_exception__15 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_exception__16 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_exception__17 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_exception__18 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_exception__19 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_exception__2 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_exception__20 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_exception__21 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_exception__22 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_exception__23 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_exception__24 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_exception__25 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_exception__26 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_exception__27 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_exception__28 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_exception__29 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_exception__3 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_exception__30 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_exception__31 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_exception__4 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_exception__5 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_exception__6 = 1'b0;
    UUT.wrapper.uut.core.rob.rob_exception__7 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_exception__8 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_exception__9 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_head = 5'b00011;
    UUT.wrapper.uut.core.rob.rob_head_lsb = 1'b0;
    UUT.wrapper.uut.core.rob.rob_state = 2'b01;
    UUT.wrapper.uut.core.rob.rob_tail = 5'b00011;
    UUT.wrapper.uut.core.rob.rob_uop_1_0_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_0_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_0_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_0_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop_1_0_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_0_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_0_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_0_ftq_idx = 3'b010;
    UUT.wrapper.uut.core.rob.rob_uop_1_0_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_0_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_0_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_0_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_0_is_rvc = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_0_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_0_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_0_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_0_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_0_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_0_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_0_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_0_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_0_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_0_uopc = 7'b1101010;
    UUT.wrapper.uut.core.rob.rob_uop_1_0_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_0_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_10_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_10_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_10_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_10_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop_1_10_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_10_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_10_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_10_ftq_idx = 3'b111;
    UUT.wrapper.uut.core.rob.rob_uop_1_10_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_10_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_10_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_10_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_10_is_rvc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_10_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_10_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_10_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_10_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_10_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_10_pc_lob = 6'b111111;
    UUT.wrapper.uut.core.rob.rob_uop_1_10_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_10_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_10_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_10_uopc = 7'b1111111;
    UUT.wrapper.uut.core.rob.rob_uop_1_10_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_10_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_11_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_11_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_11_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_11_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop_1_11_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_11_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_11_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_11_ftq_idx = 3'b111;
    UUT.wrapper.uut.core.rob.rob_uop_1_11_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_11_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_11_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_11_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_11_is_rvc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_11_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_11_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_11_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_11_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_11_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_11_pc_lob = 6'b111111;
    UUT.wrapper.uut.core.rob.rob_uop_1_11_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_11_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_11_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_11_uopc = 7'b1111111;
    UUT.wrapper.uut.core.rob.rob_uop_1_11_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_11_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_12_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_12_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_12_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_12_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop_1_12_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_12_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_12_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_12_ftq_idx = 3'b111;
    UUT.wrapper.uut.core.rob.rob_uop_1_12_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_12_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_12_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_12_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_12_is_rvc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_12_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_12_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_12_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_12_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_12_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_12_pc_lob = 6'b111111;
    UUT.wrapper.uut.core.rob.rob_uop_1_12_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_12_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_12_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_12_uopc = 7'b1111111;
    UUT.wrapper.uut.core.rob.rob_uop_1_12_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_12_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_13_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_13_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_13_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_13_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop_1_13_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_13_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_13_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_13_ftq_idx = 3'b111;
    UUT.wrapper.uut.core.rob.rob_uop_1_13_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_13_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_13_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_13_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_13_is_rvc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_13_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_13_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_13_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_13_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_13_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_13_pc_lob = 6'b111111;
    UUT.wrapper.uut.core.rob.rob_uop_1_13_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_13_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_13_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_13_uopc = 7'b1111111;
    UUT.wrapper.uut.core.rob.rob_uop_1_13_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_13_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_14_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_14_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_14_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_14_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop_1_14_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_14_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_14_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_14_ftq_idx = 3'b111;
    UUT.wrapper.uut.core.rob.rob_uop_1_14_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_14_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_14_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_14_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_14_is_rvc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_14_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_14_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_14_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_14_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_14_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_14_pc_lob = 6'b111111;
    UUT.wrapper.uut.core.rob.rob_uop_1_14_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_14_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_14_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_14_uopc = 7'b1111111;
    UUT.wrapper.uut.core.rob.rob_uop_1_14_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_14_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_15_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_15_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_15_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_15_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop_1_15_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_15_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_15_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_15_ftq_idx = 3'b111;
    UUT.wrapper.uut.core.rob.rob_uop_1_15_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_15_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_15_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_15_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_15_is_rvc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_15_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_15_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_15_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_15_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_15_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_15_pc_lob = 6'b111111;
    UUT.wrapper.uut.core.rob.rob_uop_1_15_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_15_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_15_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_15_uopc = 7'b1111111;
    UUT.wrapper.uut.core.rob.rob_uop_1_15_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_15_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_16_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_16_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_16_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_16_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop_1_16_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_16_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_16_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_16_ftq_idx = 3'b010;
    UUT.wrapper.uut.core.rob.rob_uop_1_16_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_16_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_16_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_16_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_16_is_rvc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_16_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_16_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_16_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_16_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_16_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_16_pc_lob = 6'b010000;
    UUT.wrapper.uut.core.rob.rob_uop_1_16_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_16_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_16_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_16_uopc = 7'b1101010;
    UUT.wrapper.uut.core.rob.rob_uop_1_16_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_16_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_17_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_17_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_17_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_17_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop_1_17_edge_inst = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_17_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_17_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_17_ftq_idx = 3'b000;
    UUT.wrapper.uut.core.rob.rob_uop_1_17_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_17_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_17_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_17_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_17_is_rvc = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_17_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_17_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_17_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_17_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_17_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_17_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_17_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_17_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_17_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_17_uopc = 7'b1101010;
    UUT.wrapper.uut.core.rob.rob_uop_1_17_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_17_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_18_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_18_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_18_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_18_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop_1_18_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_18_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_18_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_18_ftq_idx = 3'b111;
    UUT.wrapper.uut.core.rob.rob_uop_1_18_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_18_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_18_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_18_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_18_is_rvc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_18_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_18_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_18_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_18_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_18_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_18_pc_lob = 6'b111111;
    UUT.wrapper.uut.core.rob.rob_uop_1_18_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_18_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_18_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_18_uopc = 7'b1111111;
    UUT.wrapper.uut.core.rob.rob_uop_1_18_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_18_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_19_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_19_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_19_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_19_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop_1_19_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_19_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_19_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_19_ftq_idx = 3'b000;
    UUT.wrapper.uut.core.rob.rob_uop_1_19_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_19_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_19_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_19_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_19_is_rvc = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_19_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_19_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_19_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_19_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_19_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_19_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_19_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_19_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_19_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_19_uopc = 7'b1101010;
    UUT.wrapper.uut.core.rob.rob_uop_1_19_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_19_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_1_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_1_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_1_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_1_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop_1_1_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_1_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_1_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_1_ftq_idx = 3'b010;
    UUT.wrapper.uut.core.rob.rob_uop_1_1_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_1_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_1_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_1_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_1_is_rvc = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_1_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_1_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_1_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_1_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_1_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_1_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_1_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_1_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_1_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_1_uopc = 7'b1101010;
    UUT.wrapper.uut.core.rob.rob_uop_1_1_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_1_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_20_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_20_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_20_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_20_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop_1_20_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_20_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_20_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_20_ftq_idx = 3'b111;
    UUT.wrapper.uut.core.rob.rob_uop_1_20_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_20_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_20_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_20_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_20_is_rvc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_20_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_20_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_20_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_20_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_20_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_20_pc_lob = 6'b111111;
    UUT.wrapper.uut.core.rob.rob_uop_1_20_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_20_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_20_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_20_uopc = 7'b1111111;
    UUT.wrapper.uut.core.rob.rob_uop_1_20_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_20_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_21_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_21_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_21_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_21_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop_1_21_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_21_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_21_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_21_ftq_idx = 3'b111;
    UUT.wrapper.uut.core.rob.rob_uop_1_21_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_21_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_21_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_21_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_21_is_rvc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_21_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_21_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_21_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_21_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_21_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_21_pc_lob = 6'b111111;
    UUT.wrapper.uut.core.rob.rob_uop_1_21_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_21_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_21_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_21_uopc = 7'b1111111;
    UUT.wrapper.uut.core.rob.rob_uop_1_21_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_21_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_22_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_22_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_22_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_22_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop_1_22_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_22_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_22_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_22_ftq_idx = 3'b111;
    UUT.wrapper.uut.core.rob.rob_uop_1_22_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_22_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_22_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_22_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_22_is_rvc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_22_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_22_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_22_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_22_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_22_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_22_pc_lob = 6'b111111;
    UUT.wrapper.uut.core.rob.rob_uop_1_22_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_22_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_22_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_22_uopc = 7'b1111111;
    UUT.wrapper.uut.core.rob.rob_uop_1_22_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_22_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_23_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_23_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_23_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_23_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop_1_23_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_23_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_23_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_23_ftq_idx = 3'b111;
    UUT.wrapper.uut.core.rob.rob_uop_1_23_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_23_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_23_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_23_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_23_is_rvc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_23_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_23_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_23_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_23_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_23_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_23_pc_lob = 6'b111111;
    UUT.wrapper.uut.core.rob.rob_uop_1_23_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_23_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_23_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_23_uopc = 7'b1111111;
    UUT.wrapper.uut.core.rob.rob_uop_1_23_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_23_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_24_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_24_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_24_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_24_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop_1_24_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_24_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_24_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_24_ftq_idx = 3'b000;
    UUT.wrapper.uut.core.rob.rob_uop_1_24_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_24_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_24_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_24_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_24_is_rvc = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_24_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_24_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_24_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_24_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_24_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_24_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_24_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_24_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_24_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_24_uopc = 7'b1101010;
    UUT.wrapper.uut.core.rob.rob_uop_1_24_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_24_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_25_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_25_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_25_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_25_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop_1_25_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_25_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_25_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_25_ftq_idx = 3'b111;
    UUT.wrapper.uut.core.rob.rob_uop_1_25_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_25_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_25_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_25_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_25_is_rvc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_25_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_25_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_25_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_25_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_25_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_25_pc_lob = 6'b111111;
    UUT.wrapper.uut.core.rob.rob_uop_1_25_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_25_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_25_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_25_uopc = 7'b1111111;
    UUT.wrapper.uut.core.rob.rob_uop_1_25_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_25_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_26_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_26_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_26_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_26_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop_1_26_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_26_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_26_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_26_ftq_idx = 3'b111;
    UUT.wrapper.uut.core.rob.rob_uop_1_26_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_26_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_26_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_26_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_26_is_rvc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_26_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_26_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_26_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_26_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_26_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_26_pc_lob = 6'b111111;
    UUT.wrapper.uut.core.rob.rob_uop_1_26_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_26_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_26_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_26_uopc = 7'b1111111;
    UUT.wrapper.uut.core.rob.rob_uop_1_26_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_26_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_27_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_27_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_27_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_27_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop_1_27_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_27_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_27_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_27_ftq_idx = 3'b001;
    UUT.wrapper.uut.core.rob.rob_uop_1_27_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_27_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_27_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_27_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_27_is_rvc = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_27_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_27_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_27_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_27_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_27_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_27_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_27_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_27_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_27_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_27_uopc = 7'b1101010;
    UUT.wrapper.uut.core.rob.rob_uop_1_27_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_27_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_28_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_28_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_28_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_28_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop_1_28_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_28_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_28_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_28_ftq_idx = 3'b001;
    UUT.wrapper.uut.core.rob.rob_uop_1_28_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_28_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_28_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_28_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_28_is_rvc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_28_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_28_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_28_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_28_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_28_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_28_pc_lob = 6'b010000;
    UUT.wrapper.uut.core.rob.rob_uop_1_28_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_28_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_28_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_28_uopc = 7'b1101010;
    UUT.wrapper.uut.core.rob.rob_uop_1_28_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_28_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_29_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_29_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_29_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_29_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop_1_29_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_29_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_29_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_29_ftq_idx = 3'b010;
    UUT.wrapper.uut.core.rob.rob_uop_1_29_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_29_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_29_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_29_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_29_is_rvc = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_29_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_29_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_29_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_29_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_29_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_29_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_29_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_29_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_29_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_29_uopc = 7'b1101010;
    UUT.wrapper.uut.core.rob.rob_uop_1_29_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_29_uses_stq = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_2_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_2_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_2_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_2_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop_1_2_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_2_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_2_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_2_ftq_idx = 3'b011;
    UUT.wrapper.uut.core.rob.rob_uop_1_2_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_2_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_2_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_2_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_2_is_rvc = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_2_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_2_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_2_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_2_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_2_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_2_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_2_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_2_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_2_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_2_uopc = 7'b1101010;
    UUT.wrapper.uut.core.rob.rob_uop_1_2_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_2_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_30_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_30_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_30_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_30_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop_1_30_edge_inst = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_30_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_30_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_30_ftq_idx = 3'b101;
    UUT.wrapper.uut.core.rob.rob_uop_1_30_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_30_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_30_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_30_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_30_is_rvc = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_30_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_30_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_30_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_30_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_30_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_30_pc_lob = 6'b001100;
    UUT.wrapper.uut.core.rob.rob_uop_1_30_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_30_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_30_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_30_uopc = 7'b1101010;
    UUT.wrapper.uut.core.rob.rob_uop_1_30_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_30_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_31_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_31_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_31_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_31_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop_1_31_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_31_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_31_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_31_ftq_idx = 3'b100;
    UUT.wrapper.uut.core.rob.rob_uop_1_31_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_31_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_31_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_31_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_31_is_rvc = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_31_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_31_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_31_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_31_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_31_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_31_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_31_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_31_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_31_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_31_uopc = 7'b1101010;
    UUT.wrapper.uut.core.rob.rob_uop_1_31_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_31_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_3_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_3_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_3_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_3_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop_1_3_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_3_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_3_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_3_ftq_idx = 3'b010;
    UUT.wrapper.uut.core.rob.rob_uop_1_3_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_3_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_3_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_3_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_3_is_rvc = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_3_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_3_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_3_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_3_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_3_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_3_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_3_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_3_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_3_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_3_uopc = 7'b1101010;
    UUT.wrapper.uut.core.rob.rob_uop_1_3_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_3_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_4_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_4_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_4_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_4_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop_1_4_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_4_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_4_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_4_ftq_idx = 3'b010;
    UUT.wrapper.uut.core.rob.rob_uop_1_4_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_4_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_4_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_4_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_4_is_rvc = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_4_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_4_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_4_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_4_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_4_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_4_pc_lob = 6'b111110;
    UUT.wrapper.uut.core.rob.rob_uop_1_4_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_4_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_4_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_4_uopc = 7'b1101010;
    UUT.wrapper.uut.core.rob.rob_uop_1_4_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_4_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_5_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_5_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_5_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_5_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop_1_5_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_5_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_5_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_5_ftq_idx = 3'b111;
    UUT.wrapper.uut.core.rob.rob_uop_1_5_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_5_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_5_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_5_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_5_is_rvc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_5_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_5_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_5_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_5_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_5_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_5_pc_lob = 6'b111111;
    UUT.wrapper.uut.core.rob.rob_uop_1_5_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_5_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_5_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_5_uopc = 7'b1111111;
    UUT.wrapper.uut.core.rob.rob_uop_1_5_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_5_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_6_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_6_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_6_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_6_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop_1_6_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_6_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_6_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_6_ftq_idx = 3'b101;
    UUT.wrapper.uut.core.rob.rob_uop_1_6_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_6_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_6_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_6_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_6_is_rvc = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_6_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_6_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_6_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_6_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_6_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_6_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_6_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_6_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_6_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_6_uopc = 7'b1101010;
    UUT.wrapper.uut.core.rob.rob_uop_1_6_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_6_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_7_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_7_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_7_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_7_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop_1_7_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_7_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_7_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_7_ftq_idx = 3'b111;
    UUT.wrapper.uut.core.rob.rob_uop_1_7_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_7_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_7_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_7_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_7_is_rvc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_7_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_7_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_7_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_7_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_7_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_7_pc_lob = 6'b111111;
    UUT.wrapper.uut.core.rob.rob_uop_1_7_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_7_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_7_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_7_uopc = 7'b1111111;
    UUT.wrapper.uut.core.rob.rob_uop_1_7_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_7_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_8_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_8_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_8_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_8_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop_1_8_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_8_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_8_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_8_ftq_idx = 3'b111;
    UUT.wrapper.uut.core.rob.rob_uop_1_8_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_8_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_8_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_8_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_8_is_rvc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_8_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_8_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_8_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_8_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_8_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_8_pc_lob = 6'b111111;
    UUT.wrapper.uut.core.rob.rob_uop_1_8_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_8_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_8_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_8_uopc = 7'b1111111;
    UUT.wrapper.uut.core.rob.rob_uop_1_8_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_8_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_9_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_9_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_9_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_9_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop_1_9_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_9_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_9_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_9_ftq_idx = 3'b111;
    UUT.wrapper.uut.core.rob.rob_uop_1_9_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_9_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_9_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_9_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_9_is_rvc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_9_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_9_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_9_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop_1_9_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_9_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop_1_9_pc_lob = 6'b111111;
    UUT.wrapper.uut.core.rob.rob_uop_1_9_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_9_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_9_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop_1_9_uopc = 7'b1111111;
    UUT.wrapper.uut.core.rob.rob_uop_1_9_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop_1_9_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__0_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__0_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__0_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__0_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop__0_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__0_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__0_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__0_ftq_idx = 3'b000;
    UUT.wrapper.uut.core.rob.rob_uop__0_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__0_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__0_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__0_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__0_is_rvc = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__0_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__0_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__0_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__0_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__0_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__0_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop__0_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__0_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop__0_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__0_uopc = 7'b1101010;
    UUT.wrapper.uut.core.rob.rob_uop__0_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__0_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__10_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__10_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__10_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__10_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop__10_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__10_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__10_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__10_ftq_idx = 3'b111;
    UUT.wrapper.uut.core.rob.rob_uop__10_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__10_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__10_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__10_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__10_is_rvc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__10_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__10_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__10_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__10_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__10_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__10_pc_lob = 6'b111111;
    UUT.wrapper.uut.core.rob.rob_uop__10_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__10_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop__10_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__10_uopc = 7'b1111111;
    UUT.wrapper.uut.core.rob.rob_uop__10_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__10_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__11_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__11_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__11_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__11_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop__11_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__11_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__11_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__11_ftq_idx = 3'b111;
    UUT.wrapper.uut.core.rob.rob_uop__11_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__11_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__11_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__11_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__11_is_rvc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__11_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__11_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__11_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__11_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__11_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__11_pc_lob = 6'b111111;
    UUT.wrapper.uut.core.rob.rob_uop__11_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__11_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop__11_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__11_uopc = 7'b1111111;
    UUT.wrapper.uut.core.rob.rob_uop__11_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__11_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__12_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__12_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__12_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__12_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop__12_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__12_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__12_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__12_ftq_idx = 3'b111;
    UUT.wrapper.uut.core.rob.rob_uop__12_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__12_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__12_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__12_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__12_is_rvc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__12_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__12_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__12_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__12_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__12_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__12_pc_lob = 6'b111111;
    UUT.wrapper.uut.core.rob.rob_uop__12_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__12_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop__12_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__12_uopc = 7'b1111111;
    UUT.wrapper.uut.core.rob.rob_uop__12_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__12_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__13_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__13_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__13_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__13_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop__13_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__13_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__13_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__13_ftq_idx = 3'b111;
    UUT.wrapper.uut.core.rob.rob_uop__13_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__13_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__13_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__13_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__13_is_rvc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__13_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__13_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__13_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__13_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__13_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__13_pc_lob = 6'b111111;
    UUT.wrapper.uut.core.rob.rob_uop__13_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__13_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop__13_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__13_uopc = 7'b1111111;
    UUT.wrapper.uut.core.rob.rob_uop__13_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__13_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__14_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__14_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__14_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__14_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop__14_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__14_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__14_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__14_ftq_idx = 3'b111;
    UUT.wrapper.uut.core.rob.rob_uop__14_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__14_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__14_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__14_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__14_is_rvc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__14_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__14_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__14_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__14_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__14_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__14_pc_lob = 6'b111111;
    UUT.wrapper.uut.core.rob.rob_uop__14_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__14_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop__14_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__14_uopc = 7'b1111111;
    UUT.wrapper.uut.core.rob.rob_uop__14_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__14_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__15_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__15_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__15_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__15_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop__15_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__15_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__15_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__15_ftq_idx = 3'b111;
    UUT.wrapper.uut.core.rob.rob_uop__15_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__15_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__15_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__15_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__15_is_rvc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__15_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__15_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__15_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__15_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__15_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__15_pc_lob = 6'b111111;
    UUT.wrapper.uut.core.rob.rob_uop__15_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__15_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop__15_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__15_uopc = 7'b1111111;
    UUT.wrapper.uut.core.rob.rob_uop__15_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__15_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__16_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__16_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__16_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__16_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop__16_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__16_flush_on_commit = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__16_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__16_ftq_idx = 3'b110;
    UUT.wrapper.uut.core.rob.rob_uop__16_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__16_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__16_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__16_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__16_is_rvc = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__16_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__16_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__16_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__16_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__16_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__16_pc_lob = 6'b000100;
    UUT.wrapper.uut.core.rob.rob_uop__16_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__16_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop__16_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__16_uopc = 7'b1101010;
    UUT.wrapper.uut.core.rob.rob_uop__16_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__16_uses_stq = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__17_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__17_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__17_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__17_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop__17_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__17_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__17_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__17_ftq_idx = 3'b000;
    UUT.wrapper.uut.core.rob.rob_uop__17_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__17_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__17_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__17_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__17_is_rvc = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__17_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__17_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__17_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__17_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__17_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__17_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop__17_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__17_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop__17_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__17_uopc = 7'b0101010;
    UUT.wrapper.uut.core.rob.rob_uop__17_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__17_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__18_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__18_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__18_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__18_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop__18_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__18_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__18_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__18_ftq_idx = 3'b111;
    UUT.wrapper.uut.core.rob.rob_uop__18_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__18_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__18_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__18_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__18_is_rvc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__18_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__18_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__18_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__18_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__18_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__18_pc_lob = 6'b111111;
    UUT.wrapper.uut.core.rob.rob_uop__18_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__18_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop__18_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__18_uopc = 7'b1111111;
    UUT.wrapper.uut.core.rob.rob_uop__18_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__18_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__19_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__19_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__19_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__19_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop__19_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__19_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__19_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__19_ftq_idx = 3'b000;
    UUT.wrapper.uut.core.rob.rob_uop__19_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__19_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__19_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__19_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__19_is_rvc = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__19_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__19_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__19_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__19_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__19_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__19_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop__19_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__19_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop__19_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__19_uopc = 7'b0101010;
    UUT.wrapper.uut.core.rob.rob_uop__19_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__19_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__1_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__1_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__1_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__1_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop__1_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__1_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__1_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__1_ftq_idx = 3'b000;
    UUT.wrapper.uut.core.rob.rob_uop__1_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__1_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__1_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__1_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__1_is_rvc = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__1_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__1_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__1_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__1_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__1_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__1_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop__1_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__1_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop__1_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__1_uopc = 7'b1101010;
    UUT.wrapper.uut.core.rob.rob_uop__1_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__1_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__20_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__20_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__20_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__20_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop__20_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__20_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__20_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__20_ftq_idx = 3'b111;
    UUT.wrapper.uut.core.rob.rob_uop__20_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__20_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__20_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__20_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__20_is_rvc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__20_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__20_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__20_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__20_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__20_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__20_pc_lob = 6'b111111;
    UUT.wrapper.uut.core.rob.rob_uop__20_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__20_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop__20_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__20_uopc = 7'b1111111;
    UUT.wrapper.uut.core.rob.rob_uop__20_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__20_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__21_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__21_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__21_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__21_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop__21_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__21_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__21_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__21_ftq_idx = 3'b111;
    UUT.wrapper.uut.core.rob.rob_uop__21_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__21_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__21_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__21_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__21_is_rvc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__21_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__21_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__21_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__21_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__21_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__21_pc_lob = 6'b111111;
    UUT.wrapper.uut.core.rob.rob_uop__21_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__21_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop__21_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__21_uopc = 7'b1111111;
    UUT.wrapper.uut.core.rob.rob_uop__21_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__21_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__22_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__22_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__22_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__22_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop__22_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__22_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__22_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__22_ftq_idx = 3'b111;
    UUT.wrapper.uut.core.rob.rob_uop__22_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__22_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__22_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__22_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__22_is_rvc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__22_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__22_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__22_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__22_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__22_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__22_pc_lob = 6'b111111;
    UUT.wrapper.uut.core.rob.rob_uop__22_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__22_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop__22_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__22_uopc = 7'b1111111;
    UUT.wrapper.uut.core.rob.rob_uop__22_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__22_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__23_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__23_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__23_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__23_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop__23_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__23_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__23_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__23_ftq_idx = 3'b111;
    UUT.wrapper.uut.core.rob.rob_uop__23_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__23_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__23_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__23_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__23_is_rvc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__23_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__23_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__23_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__23_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__23_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__23_pc_lob = 6'b111111;
    UUT.wrapper.uut.core.rob.rob_uop__23_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__23_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop__23_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__23_uopc = 7'b1111111;
    UUT.wrapper.uut.core.rob.rob_uop__23_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__23_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__24_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__24_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__24_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__24_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop__24_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__24_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__24_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__24_ftq_idx = 3'b000;
    UUT.wrapper.uut.core.rob.rob_uop__24_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__24_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__24_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__24_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__24_is_rvc = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__24_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__24_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__24_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__24_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__24_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__24_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop__24_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__24_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop__24_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__24_uopc = 7'b0101010;
    UUT.wrapper.uut.core.rob.rob_uop__24_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__24_uses_stq = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__25_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__25_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__25_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__25_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop__25_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__25_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__25_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__25_ftq_idx = 3'b111;
    UUT.wrapper.uut.core.rob.rob_uop__25_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__25_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__25_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__25_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__25_is_rvc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__25_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__25_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__25_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__25_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__25_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__25_pc_lob = 6'b111111;
    UUT.wrapper.uut.core.rob.rob_uop__25_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__25_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop__25_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__25_uopc = 7'b1111111;
    UUT.wrapper.uut.core.rob.rob_uop__25_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__25_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__26_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__26_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__26_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__26_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop__26_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__26_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__26_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__26_ftq_idx = 3'b111;
    UUT.wrapper.uut.core.rob.rob_uop__26_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__26_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__26_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__26_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__26_is_rvc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__26_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__26_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__26_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__26_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__26_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__26_pc_lob = 6'b111111;
    UUT.wrapper.uut.core.rob.rob_uop__26_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__26_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop__26_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__26_uopc = 7'b1111111;
    UUT.wrapper.uut.core.rob.rob_uop__26_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__26_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__27_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__27_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__27_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__27_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop__27_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__27_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__27_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__27_ftq_idx = 3'b000;
    UUT.wrapper.uut.core.rob.rob_uop__27_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__27_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__27_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__27_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__27_is_rvc = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__27_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__27_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__27_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__27_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__27_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__27_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop__27_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__27_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop__27_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__27_uopc = 7'b0101010;
    UUT.wrapper.uut.core.rob.rob_uop__27_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__27_uses_stq = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__28_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__28_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__28_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__28_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop__28_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__28_flush_on_commit = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__28_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__28_ftq_idx = 3'b110;
    UUT.wrapper.uut.core.rob.rob_uop__28_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__28_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__28_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__28_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__28_is_rvc = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__28_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__28_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__28_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__28_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__28_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__28_pc_lob = 6'b000100;
    UUT.wrapper.uut.core.rob.rob_uop__28_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__28_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop__28_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__28_uopc = 7'b1101010;
    UUT.wrapper.uut.core.rob.rob_uop__28_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__28_uses_stq = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__29_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__29_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__29_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__29_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop__29_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__29_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__29_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__29_ftq_idx = 3'b000;
    UUT.wrapper.uut.core.rob.rob_uop__29_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__29_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__29_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__29_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__29_is_rvc = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__29_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__29_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__29_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__29_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__29_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__29_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop__29_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__29_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop__29_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__29_uopc = 7'b1101010;
    UUT.wrapper.uut.core.rob.rob_uop__29_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__29_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__2_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__2_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__2_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__2_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop__2_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__2_flush_on_commit = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__2_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__2_ftq_idx = 3'b110;
    UUT.wrapper.uut.core.rob.rob_uop__2_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__2_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__2_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__2_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__2_is_rvc = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__2_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__2_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__2_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__2_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__2_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__2_pc_lob = 6'b000100;
    UUT.wrapper.uut.core.rob.rob_uop__2_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__2_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop__2_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__2_uopc = 7'b1101010;
    UUT.wrapper.uut.core.rob.rob_uop__2_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__2_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__30_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__30_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__30_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__30_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop__30_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__30_flush_on_commit = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__30_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__30_ftq_idx = 3'b110;
    UUT.wrapper.uut.core.rob.rob_uop__30_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__30_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__30_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__30_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__30_is_rvc = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__30_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__30_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__30_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__30_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__30_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__30_pc_lob = 6'b000010;
    UUT.wrapper.uut.core.rob.rob_uop__30_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__30_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop__30_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__30_uopc = 7'b1101010;
    UUT.wrapper.uut.core.rob.rob_uop__30_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__30_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__31_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__31_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__31_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__31_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop__31_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__31_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__31_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__31_ftq_idx = 3'b000;
    UUT.wrapper.uut.core.rob.rob_uop__31_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__31_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__31_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__31_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__31_is_rvc = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__31_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__31_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__31_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__31_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__31_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__31_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop__31_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__31_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop__31_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__31_uopc = 7'b1101010;
    UUT.wrapper.uut.core.rob.rob_uop__31_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__31_uses_stq = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__3_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__3_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__3_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__3_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop__3_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__3_flush_on_commit = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__3_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__3_ftq_idx = 3'b000;
    UUT.wrapper.uut.core.rob.rob_uop__3_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__3_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__3_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__3_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__3_is_rvc = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__3_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__3_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__3_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__3_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__3_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__3_pc_lob = 6'b100000;
    UUT.wrapper.uut.core.rob.rob_uop__3_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__3_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop__3_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__3_uopc = 7'b1101010;
    UUT.wrapper.uut.core.rob.rob_uop__3_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__3_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__4_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__4_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__4_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__4_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop__4_edge_inst = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__4_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__4_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__4_ftq_idx = 3'b000;
    UUT.wrapper.uut.core.rob.rob_uop__4_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__4_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__4_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__4_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__4_is_rvc = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__4_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__4_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__4_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__4_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__4_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__4_pc_lob = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop__4_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__4_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop__4_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__4_uopc = 7'b0101010;
    UUT.wrapper.uut.core.rob.rob_uop__4_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__4_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__5_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__5_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__5_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__5_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop__5_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__5_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__5_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__5_ftq_idx = 3'b111;
    UUT.wrapper.uut.core.rob.rob_uop__5_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__5_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__5_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__5_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__5_is_rvc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__5_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__5_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__5_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__5_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__5_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__5_pc_lob = 6'b111111;
    UUT.wrapper.uut.core.rob.rob_uop__5_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__5_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop__5_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__5_uopc = 7'b1111111;
    UUT.wrapper.uut.core.rob.rob_uop__5_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__5_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__6_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__6_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__6_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__6_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop__6_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__6_flush_on_commit = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__6_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__6_ftq_idx = 3'b000;
    UUT.wrapper.uut.core.rob.rob_uop__6_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__6_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__6_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__6_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__6_is_rvc = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__6_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__6_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__6_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__6_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__6_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__6_pc_lob = 6'b000100;
    UUT.wrapper.uut.core.rob.rob_uop__6_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__6_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop__6_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__6_uopc = 7'b1101010;
    UUT.wrapper.uut.core.rob.rob_uop__6_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__6_uses_stq = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__7_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__7_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__7_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__7_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop__7_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__7_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__7_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__7_ftq_idx = 3'b111;
    UUT.wrapper.uut.core.rob.rob_uop__7_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__7_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__7_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__7_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__7_is_rvc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__7_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__7_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__7_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__7_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__7_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__7_pc_lob = 6'b111111;
    UUT.wrapper.uut.core.rob.rob_uop__7_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__7_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop__7_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__7_uopc = 7'b1111111;
    UUT.wrapper.uut.core.rob.rob_uop__7_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__7_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__8_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__8_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__8_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__8_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop__8_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__8_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__8_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__8_ftq_idx = 3'b111;
    UUT.wrapper.uut.core.rob.rob_uop__8_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__8_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__8_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__8_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__8_is_rvc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__8_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__8_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__8_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__8_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__8_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__8_pc_lob = 6'b111111;
    UUT.wrapper.uut.core.rob.rob_uop__8_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__8_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop__8_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__8_uopc = 7'b1111111;
    UUT.wrapper.uut.core.rob.rob_uop__8_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__8_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__9_br_mask = 12'b000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__9_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__9_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_uop__9_dst_rtype = 2'b00;
    UUT.wrapper.uut.core.rob.rob_uop__9_edge_inst = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__9_flush_on_commit = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__9_fp_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__9_ftq_idx = 3'b111;
    UUT.wrapper.uut.core.rob.rob_uop__9_is_br = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__9_is_fencei = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__9_is_jal = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__9_is_jalr = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__9_is_rvc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__9_is_sys_pc2epc = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__9_ldst = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__9_ldst_val = 1'b0;
    UUT.wrapper.uut.core.rob.rob_uop__9_lrs1 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__9_lrs2 = 5'b00000;
    UUT.wrapper.uut.core.rob.rob_uop__9_pc_lob = 6'b111111;
    UUT.wrapper.uut.core.rob.rob_uop__9_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__9_rob_idx = 6'b000000;
    UUT.wrapper.uut.core.rob.rob_uop__9_stale_pdst = 7'b0000000;
    UUT.wrapper.uut.core.rob.rob_uop__9_uopc = 7'b1111111;
    UUT.wrapper.uut.core.rob.rob_uop__9_uses_ldq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_uop__9_uses_stq = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val_1_0 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val_1_1 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val_1_10 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val_1_11 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val_1_12 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val_1_13 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val_1_14 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val_1_15 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val_1_16 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val_1_17 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val_1_18 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val_1_19 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val_1_2 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val_1_20 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val_1_21 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val_1_22 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val_1_23 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val_1_24 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val_1_25 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val_1_26 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val_1_27 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val_1_28 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val_1_29 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val_1_3 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val_1_30 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val_1_31 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val_1_4 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val_1_5 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val_1_6 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val_1_7 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val_1_8 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val_1_9 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val__0 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val__1 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val__10 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val__11 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val__12 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val__13 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val__14 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val__15 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val__16 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val__17 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val__18 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val__19 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val__2 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val__20 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val__21 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val__22 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val__23 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val__24 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val__25 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val__26 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val__27 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val__28 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val__29 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val__3 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val__30 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val__31 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val__4 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val__5 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val__6 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val__7 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val__8 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_val__9 = 1'b1;
    UUT.wrapper.uut.core.saturating_loads_counter = 5'b11111;
    UUT.wrapper.uut.dcache.beatsLeft = 3'b111;
    UUT.wrapper.uut.dcache.data.array_0_0_0_io_resp_0_0_MPORT_addr_pipe_0 = 4'b1110;
    UUT.wrapper.uut.dcache.data.io_resp_0_0_REG = 64'b0000000000000000101000000000000010101000000000000000000000000001;
    UUT.wrapper.uut.dcache.io_lsu_perf_acquire_counter = 3'b111;
    UUT.wrapper.uut.dcache.io_lsu_perf_release_counter = 3'b001;
    UUT.wrapper.uut.dcache.lrsc_addr = 34'b0000000000010000000000000000000000;
    UUT.wrapper.uut.dcache.lrsc_count = 7'b1111111;
    UUT.wrapper.uut.dcache.meta_0.rst_cnt = 2'b01;
    UUT.wrapper.uut.dcache.meta_0.tag_array_0_MPORT_1_addr_pipe_0 = 1'b1;
    UUT.wrapper.uut.dcache.mshrs.beatsLeft = 3'b111;
    UUT.wrapper.uut.dcache.mshrs.beatsLeft_1 = 1'b0;
    UUT.wrapper.uut.dcache.mshrs.mmios_0.grant_word = 64'b1111111111111111111111111111111111111111111111101000000000000000;
    UUT.wrapper.uut.dcache.mshrs.mmios_0.req_addr = 40'b1111111111111111111111111111111111111000;
    UUT.wrapper.uut.dcache.mshrs.mmios_0.req_data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.dcache.mshrs.mmios_0.req_is_hella = 1'b1;
    UUT.wrapper.uut.dcache.mshrs.mmios_0.req_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.dcache.mshrs.mmios_0.req_uop_is_amo = 1'b0;
    UUT.wrapper.uut.dcache.mshrs.mmios_0.req_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.dcache.mshrs.mmios_0.req_uop_mem_cmd = 5'b11111;
    UUT.wrapper.uut.dcache.mshrs.mmios_0.req_uop_mem_signed = 1'b1;
    UUT.wrapper.uut.dcache.mshrs.mmios_0.req_uop_mem_size = 2'b11;
    UUT.wrapper.uut.dcache.mshrs.mmios_0.req_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.dcache.mshrs.mmios_0.req_uop_uses_ldq = 1'b0;
    UUT.wrapper.uut.dcache.mshrs.mmios_0.req_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.dcache.mshrs.mmios_0.state = 2'b00;
    UUT.wrapper.uut.dcache.mshrs.mshr_alloc_idx_REG = 1'b0;
    UUT.wrapper.uut.dcache.mshrs.mshr_head = 1'b0;
    UUT.wrapper.uut.dcache.mshrs.mshrs_0.commit_line = 1'b0;
    UUT.wrapper.uut.dcache.mshrs.mshrs_0.counter = 3'b111;
    UUT.wrapper.uut.dcache.mshrs.mshrs_0.grant_had_data = 1'b0;
    UUT.wrapper.uut.dcache.mshrs.mshrs_0.grantack_bits_sink = 2'b00;
    UUT.wrapper.uut.dcache.mshrs.mshrs_0.grantack_valid = 1'b0;
    UUT.wrapper.uut.dcache.mshrs.mshrs_0.meta_hazard = 2'b00;
    UUT.wrapper.uut.dcache.mshrs.mshrs_0.new_coh_state = 2'b00;
    UUT.wrapper.uut.dcache.mshrs.mshrs_0.refill_ctr = 3'b000;
    UUT.wrapper.uut.dcache.mshrs.mshrs_0.req_addr = 40'b1000000011111111111111111111111111111111;
    UUT.wrapper.uut.dcache.mshrs.mshrs_0.req_old_meta_coh_state = 2'b00;
    UUT.wrapper.uut.dcache.mshrs.mshrs_0.req_old_meta_tag = 25'b0000000000000000000000000;
    UUT.wrapper.uut.dcache.mshrs.mshrs_0.req_uop_mem_cmd = 5'b10001;
    UUT.wrapper.uut.dcache.mshrs.mshrs_0.req_way_en = 1'b1;
    UUT.wrapper.uut.dcache.mshrs.mshrs_0.rpq.deq_ptr_value = 1'b1;
    UUT.wrapper.uut.dcache.mshrs.mshrs_0.rpq.enq_ptr_value = 1'b1;
    UUT.wrapper.uut.dcache.mshrs.mshrs_0.rpq.maybe_full = 1'b1;
    UUT.wrapper.uut.dcache.mshrs.mshrs_0.rpq.uops_0_br_mask = 12'b111111111111;
    UUT.wrapper.uut.dcache.mshrs.mshrs_0.rpq.uops_0_is_amo = 1'b0;
    UUT.wrapper.uut.dcache.mshrs.mshrs_0.rpq.uops_0_ldq_idx = 4'b0000;
    UUT.wrapper.uut.dcache.mshrs.mshrs_0.rpq.uops_0_mem_cmd = 5'b00000;
    UUT.wrapper.uut.dcache.mshrs.mshrs_0.rpq.uops_0_mem_signed = 1'b0;
    UUT.wrapper.uut.dcache.mshrs.mshrs_0.rpq.uops_0_mem_size = 2'b00;
    UUT.wrapper.uut.dcache.mshrs.mshrs_0.rpq.uops_0_stq_idx = 4'b0000;
    UUT.wrapper.uut.dcache.mshrs.mshrs_0.rpq.uops_0_uses_ldq = 1'b0;
    UUT.wrapper.uut.dcache.mshrs.mshrs_0.rpq.uops_0_uses_stq = 1'b0;
    UUT.wrapper.uut.dcache.mshrs.mshrs_0.rpq.uops_1_br_mask = 12'b111111111111;
    UUT.wrapper.uut.dcache.mshrs.mshrs_0.rpq.uops_1_is_amo = 1'b0;
    UUT.wrapper.uut.dcache.mshrs.mshrs_0.rpq.uops_1_ldq_idx = 4'b0000;
    UUT.wrapper.uut.dcache.mshrs.mshrs_0.rpq.uops_1_mem_cmd = 5'b00000;
    UUT.wrapper.uut.dcache.mshrs.mshrs_0.rpq.uops_1_mem_signed = 1'b0;
    UUT.wrapper.uut.dcache.mshrs.mshrs_0.rpq.uops_1_mem_size = 2'b00;
    UUT.wrapper.uut.dcache.mshrs.mshrs_0.rpq.uops_1_stq_idx = 4'b0000;
    UUT.wrapper.uut.dcache.mshrs.mshrs_0.rpq.uops_1_uses_ldq = 1'b0;
    UUT.wrapper.uut.dcache.mshrs.mshrs_0.rpq.uops_1_uses_stq = 1'b0;
    UUT.wrapper.uut.dcache.mshrs.mshrs_0.rpq.valids_0 = 1'b0;
    UUT.wrapper.uut.dcache.mshrs.mshrs_0.rpq.valids_1 = 1'b1;
    UUT.wrapper.uut.dcache.mshrs.mshrs_0.state = 5'b11111;
    UUT.wrapper.uut.dcache.mshrs.mshrs_1.commit_line = 1'b0;
    UUT.wrapper.uut.dcache.mshrs.mshrs_1.counter = 3'b111;
    UUT.wrapper.uut.dcache.mshrs.mshrs_1.grant_had_data = 1'b0;
    UUT.wrapper.uut.dcache.mshrs.mshrs_1.grantack_bits_sink = 2'b00;
    UUT.wrapper.uut.dcache.mshrs.mshrs_1.grantack_valid = 1'b0;
    UUT.wrapper.uut.dcache.mshrs.mshrs_1.meta_hazard = 2'b00;
    UUT.wrapper.uut.dcache.mshrs.mshrs_1.new_coh_state = 2'b00;
    UUT.wrapper.uut.dcache.mshrs.mshrs_1.refill_ctr = 3'b000;
    UUT.wrapper.uut.dcache.mshrs.mshrs_1.req_addr = 40'b0000000011111111111111111111111111111111;
    UUT.wrapper.uut.dcache.mshrs.mshrs_1.req_old_meta_coh_state = 2'b00;
    UUT.wrapper.uut.dcache.mshrs.mshrs_1.req_old_meta_tag = 25'b0000000000000000000000000;
    UUT.wrapper.uut.dcache.mshrs.mshrs_1.req_uop_mem_cmd = 5'b10001;
    UUT.wrapper.uut.dcache.mshrs.mshrs_1.req_way_en = 1'b1;
    UUT.wrapper.uut.dcache.mshrs.mshrs_1.rpq.deq_ptr_value = 1'b1;
    UUT.wrapper.uut.dcache.mshrs.mshrs_1.rpq.enq_ptr_value = 1'b1;
    UUT.wrapper.uut.dcache.mshrs.mshrs_1.rpq.maybe_full = 1'b1;
    UUT.wrapper.uut.dcache.mshrs.mshrs_1.rpq.uops_0_br_mask = 12'b111111111111;
    UUT.wrapper.uut.dcache.mshrs.mshrs_1.rpq.uops_0_is_amo = 1'b0;
    UUT.wrapper.uut.dcache.mshrs.mshrs_1.rpq.uops_0_ldq_idx = 4'b0000;
    UUT.wrapper.uut.dcache.mshrs.mshrs_1.rpq.uops_0_mem_cmd = 5'b00000;
    UUT.wrapper.uut.dcache.mshrs.mshrs_1.rpq.uops_0_mem_signed = 1'b0;
    UUT.wrapper.uut.dcache.mshrs.mshrs_1.rpq.uops_0_mem_size = 2'b00;
    UUT.wrapper.uut.dcache.mshrs.mshrs_1.rpq.uops_0_stq_idx = 4'b0000;
    UUT.wrapper.uut.dcache.mshrs.mshrs_1.rpq.uops_0_uses_ldq = 1'b0;
    UUT.wrapper.uut.dcache.mshrs.mshrs_1.rpq.uops_0_uses_stq = 1'b0;
    UUT.wrapper.uut.dcache.mshrs.mshrs_1.rpq.uops_1_br_mask = 12'b111111111111;
    UUT.wrapper.uut.dcache.mshrs.mshrs_1.rpq.uops_1_is_amo = 1'b0;
    UUT.wrapper.uut.dcache.mshrs.mshrs_1.rpq.uops_1_ldq_idx = 4'b0000;
    UUT.wrapper.uut.dcache.mshrs.mshrs_1.rpq.uops_1_mem_cmd = 5'b00000;
    UUT.wrapper.uut.dcache.mshrs.mshrs_1.rpq.uops_1_mem_signed = 1'b0;
    UUT.wrapper.uut.dcache.mshrs.mshrs_1.rpq.uops_1_mem_size = 2'b00;
    UUT.wrapper.uut.dcache.mshrs.mshrs_1.rpq.uops_1_stq_idx = 4'b0000;
    UUT.wrapper.uut.dcache.mshrs.mshrs_1.rpq.uops_1_uses_ldq = 1'b0;
    UUT.wrapper.uut.dcache.mshrs.mshrs_1.rpq.uops_1_uses_stq = 1'b0;
    UUT.wrapper.uut.dcache.mshrs.mshrs_1.rpq.valids_0 = 1'b1;
    UUT.wrapper.uut.dcache.mshrs.mshrs_1.rpq.valids_1 = 1'b1;
    UUT.wrapper.uut.dcache.mshrs.mshrs_1.state = 5'b00001;
    UUT.wrapper.uut.dcache.mshrs.respq.deq_ptr_value = 2'b11;
    UUT.wrapper.uut.dcache.mshrs.respq.enq_ptr_value = 2'b11;
    UUT.wrapper.uut.dcache.mshrs.respq.maybe_full = 1'b1;
    UUT.wrapper.uut.dcache.mshrs.respq.uops_0_br_mask = 12'b111111111111;
    UUT.wrapper.uut.dcache.mshrs.respq.uops_0_is_amo = 1'b1;
    UUT.wrapper.uut.dcache.mshrs.respq.uops_0_ldq_idx = 4'b1111;
    UUT.wrapper.uut.dcache.mshrs.respq.uops_0_stq_idx = 4'b1111;
    UUT.wrapper.uut.dcache.mshrs.respq.uops_0_uses_ldq = 1'b1;
    UUT.wrapper.uut.dcache.mshrs.respq.uops_0_uses_stq = 1'b1;
    UUT.wrapper.uut.dcache.mshrs.respq.uops_1_br_mask = 12'b111111111111;
    UUT.wrapper.uut.dcache.mshrs.respq.uops_1_is_amo = 1'b1;
    UUT.wrapper.uut.dcache.mshrs.respq.uops_1_ldq_idx = 4'b1111;
    UUT.wrapper.uut.dcache.mshrs.respq.uops_1_stq_idx = 4'b1111;
    UUT.wrapper.uut.dcache.mshrs.respq.uops_1_uses_ldq = 1'b1;
    UUT.wrapper.uut.dcache.mshrs.respq.uops_1_uses_stq = 1'b1;
    UUT.wrapper.uut.dcache.mshrs.respq.uops_2_br_mask = 12'b111111111111;
    UUT.wrapper.uut.dcache.mshrs.respq.uops_2_is_amo = 1'b1;
    UUT.wrapper.uut.dcache.mshrs.respq.uops_2_ldq_idx = 4'b1111;
    UUT.wrapper.uut.dcache.mshrs.respq.uops_2_stq_idx = 4'b1111;
    UUT.wrapper.uut.dcache.mshrs.respq.uops_2_uses_ldq = 1'b1;
    UUT.wrapper.uut.dcache.mshrs.respq.uops_2_uses_stq = 1'b1;
    UUT.wrapper.uut.dcache.mshrs.respq.uops_3_br_mask = 12'b101011010010;
    UUT.wrapper.uut.dcache.mshrs.respq.uops_3_is_amo = 1'b1;
    UUT.wrapper.uut.dcache.mshrs.respq.uops_3_ldq_idx = 4'b0011;
    UUT.wrapper.uut.dcache.mshrs.respq.uops_3_stq_idx = 4'b0000;
    UUT.wrapper.uut.dcache.mshrs.respq.uops_3_uses_ldq = 1'b1;
    UUT.wrapper.uut.dcache.mshrs.respq.uops_3_uses_stq = 1'b1;
    UUT.wrapper.uut.dcache.mshrs.respq.valids_0 = 1'b1;
    UUT.wrapper.uut.dcache.mshrs.respq.valids_1 = 1'b1;
    UUT.wrapper.uut.dcache.mshrs.respq.valids_2 = 1'b1;
    UUT.wrapper.uut.dcache.mshrs.respq.valids_3 = 1'b1;
    UUT.wrapper.uut.dcache.mshrs.sdq_val = 2'b11;
    UUT.wrapper.uut.dcache.mshrs.state_1_0 = 1'b0;
    UUT.wrapper.uut.dcache.mshrs.state_1_1 = 1'b0;
    UUT.wrapper.uut.dcache.mshrs.state__0 = 1'b1;
    UUT.wrapper.uut.dcache.mshrs.state__1 = 1'b1;
    UUT.wrapper.uut.dcache.mshrs.state__2 = 1'b1;
    UUT.wrapper.uut.dcache.mshrs_io_meta_resp_bits_REG_0_coh_state = 2'b00;
    UUT.wrapper.uut.dcache.prober.old_coh_state = 2'b00;
    UUT.wrapper.uut.dcache.prober.req_address = 32'b00000000000000000000000000111111;
    UUT.wrapper.uut.dcache.prober.req_param = 2'b11;
    UUT.wrapper.uut.dcache.prober.req_size = 3'b111;
    UUT.wrapper.uut.dcache.prober.req_source = 2'b00;
    UUT.wrapper.uut.dcache.prober.state = 4'b0111;
    UUT.wrapper.uut.dcache.prober.way_en = 1'b1;
    UUT.wrapper.uut.dcache.s1_mshr_meta_read_way_en = 1'b1;
    UUT.wrapper.uut.dcache.s1_replay_way_en = 1'b1;
    UUT.wrapper.uut.dcache.s1_req_0_addr = 40'b0000000011111111111111101111111111111111;
    UUT.wrapper.uut.dcache.s1_req_0_data = 64'b1111111111111111111111111111111100000001000000010000000000000000;
    UUT.wrapper.uut.dcache.s1_req_0_is_hella = 1'b1;
    UUT.wrapper.uut.dcache.s1_req_0_uop_br_mask = 12'b111111111111;
    UUT.wrapper.uut.dcache.s1_req_0_uop_is_amo = 1'b1;
    UUT.wrapper.uut.dcache.s1_req_0_uop_ldq_idx = 4'b1111;
    UUT.wrapper.uut.dcache.s1_req_0_uop_mem_cmd = 5'b11111;
    UUT.wrapper.uut.dcache.s1_req_0_uop_mem_signed = 1'b1;
    UUT.wrapper.uut.dcache.s1_req_0_uop_mem_size = 2'b01;
    UUT.wrapper.uut.dcache.s1_req_0_uop_stq_idx = 4'b1111;
    UUT.wrapper.uut.dcache.s1_req_0_uop_uses_ldq = 1'b1;
    UUT.wrapper.uut.dcache.s1_req_0_uop_uses_stq = 1'b1;
    UUT.wrapper.uut.dcache.s1_send_resp_or_nack_0 = 1'b1;
    UUT.wrapper.uut.dcache.s1_type = 3'b111;
    UUT.wrapper.uut.dcache.s1_valid_REG = 1'b1;
    UUT.wrapper.uut.dcache.s1_wb_way_en = 1'b1;
    UUT.wrapper.uut.dcache.s2_hit_state_REG_state = 2'b11;
    UUT.wrapper.uut.dcache.s2_lr_REG = 1'b0;
    UUT.wrapper.uut.dcache.s2_nack_hit_0 = 1'b0;
    UUT.wrapper.uut.dcache.s2_repl_meta_REG_coh_state = 2'b00;
    UUT.wrapper.uut.dcache.s2_repl_meta_REG_tag = 25'b0000000000000000000000000;
    UUT.wrapper.uut.dcache.s2_req_0_addr = 40'b0000000011111111111111111111111111111101;
    UUT.wrapper.uut.dcache.s2_req_0_data = 64'b1011111111111111010111111111111011100101000000000000000000000001;
    UUT.wrapper.uut.dcache.s2_req_0_is_hella = 1'b1;
    UUT.wrapper.uut.dcache.s2_req_0_uop_br_mask = 12'b101011010010;
    UUT.wrapper.uut.dcache.s2_req_0_uop_is_amo = 1'b1;
    UUT.wrapper.uut.dcache.s2_req_0_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.dcache.s2_req_0_uop_mem_cmd = 5'b11111;
    UUT.wrapper.uut.dcache.s2_req_0_uop_mem_signed = 1'b0;
    UUT.wrapper.uut.dcache.s2_req_0_uop_mem_size = 2'b00;
    UUT.wrapper.uut.dcache.s2_req_0_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.dcache.s2_req_0_uop_uses_ldq = 1'b1;
    UUT.wrapper.uut.dcache.s2_req_0_uop_uses_stq = 1'b1;
    UUT.wrapper.uut.dcache.s2_sc_REG = 1'b0;
    UUT.wrapper.uut.dcache.s2_send_nack_REG = 1'b0;
    UUT.wrapper.uut.dcache.s2_send_resp_REG = 1'b0;
    UUT.wrapper.uut.dcache.s2_tag_match_way_0 = 1'b1;
    UUT.wrapper.uut.dcache.s2_type = 3'b010;
    UUT.wrapper.uut.dcache.s2_valid_REG = 1'b1;
    UUT.wrapper.uut.dcache.s2_wb_idx_matches_0 = 1'b0;
    UUT.wrapper.uut.dcache.s3_req_addr = 40'b0000000011111111111111101111111111111111;
    UUT.wrapper.uut.dcache.s3_req_data = 64'b0000000000000000000000000000000000000001000000010000000000000001;
    UUT.wrapper.uut.dcache.s3_valid = 1'b1;
    UUT.wrapper.uut.dcache.s3_way = 1'b1;
    UUT.wrapper.uut.dcache.s4_req_addr = 40'b0000000011111111111111101111111111111111;
    UUT.wrapper.uut.dcache.s4_req_data = 64'b0000000000000000000000000000000010000000000000000000000000000000;
    UUT.wrapper.uut.dcache.s4_valid = 1'b1;
    UUT.wrapper.uut.dcache.s5_req_addr = 40'b0000000011111111111111111111111111111111;
    UUT.wrapper.uut.dcache.s5_req_data = 64'b0000000000000000000000000000000010100000000000000000000010000010;
    UUT.wrapper.uut.dcache.s5_valid = 1'b0;
    UUT.wrapper.uut.dcache.state_0 = 1'b1;
    UUT.wrapper.uut.dcache.state_1 = 1'b1;
    UUT.wrapper.uut.dcache.wb.acked = 1'b0;
    UUT.wrapper.uut.dcache.wb.data_req_cnt = 4'b0000;
    UUT.wrapper.uut.dcache.wb.r1_data_req_cnt = 4'b0000;
    UUT.wrapper.uut.dcache.wb.r1_data_req_fired = 1'b0;
    UUT.wrapper.uut.dcache.wb.r2_data_req_cnt = 4'b0000;
    UUT.wrapper.uut.dcache.wb.r2_data_req_fired = 1'b0;
    UUT.wrapper.uut.dcache.wb.req_idx = 1'b1;
    UUT.wrapper.uut.dcache.wb.req_param = 3'b000;
    UUT.wrapper.uut.dcache.wb.req_tag = 25'b0000000000000000000000000;
    UUT.wrapper.uut.dcache.wb.req_voluntary = 1'b0;
    UUT.wrapper.uut.dcache.wb.req_way_en = 1'b1;
    UUT.wrapper.uut.dcache.wb.state = 3'b111;
    UUT.wrapper.uut.dcache.wb.wb_buffer_0 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.dcache.wb.wb_buffer_1 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.dcache.wb.wb_buffer_2 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.dcache.wb.wb_buffer_3 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.dcache.wb.wb_buffer_4 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.dcache.wb.wb_buffer_5 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.dcache.wb.wb_buffer_6 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.dcache.wb.wb_buffer_7 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.frontend.REG = 1'b0;
    UUT.wrapper.uut.frontend.f3.maybe_full = 1'b1;
    UUT.wrapper.uut.frontend.f3_bpd_resp.maybe_full = 1'b1;
    UUT.wrapper.uut.frontend.f3_bpd_resp_io_enq_valid_REG = 1'b0;
    UUT.wrapper.uut.frontend.f3_prev_half = 16'b1001110000000010;
    UUT.wrapper.uut.frontend.f3_prev_is_half = 1'b1;
    UUT.wrapper.uut.frontend.f4.maybe_full = 1'b1;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_0_bp_debug_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_0_bp_xcpt_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_0_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_0_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_0_edge_inst = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_0_ftq_idx = 3'b000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_0_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_0_is_rvc = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_0_is_sfb = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_0_pc_lob = 6'b000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_0_taken = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_0_xcpt_ae_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_0_xcpt_pf_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_10_bp_debug_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_10_bp_xcpt_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_10_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_10_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_10_edge_inst = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_10_ftq_idx = 3'b000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_10_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_10_is_rvc = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_10_is_sfb = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_10_pc_lob = 6'b000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_10_taken = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_10_xcpt_ae_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_10_xcpt_pf_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_11_bp_debug_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_11_bp_xcpt_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_11_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_11_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_11_edge_inst = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_11_ftq_idx = 3'b111;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_11_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_11_is_rvc = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_11_is_sfb = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_11_pc_lob = 6'b000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_11_taken = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_11_xcpt_ae_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_11_xcpt_pf_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_12_bp_debug_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_12_bp_xcpt_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_12_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_12_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_12_edge_inst = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_12_ftq_idx = 3'b000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_12_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_12_is_rvc = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_12_is_sfb = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_12_pc_lob = 6'b000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_12_taken = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_12_xcpt_ae_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_12_xcpt_pf_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_13_bp_debug_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_13_bp_xcpt_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_13_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_13_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_13_edge_inst = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_13_ftq_idx = 3'b111;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_13_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_13_is_rvc = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_13_is_sfb = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_13_pc_lob = 6'b000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_13_taken = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_13_xcpt_ae_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_13_xcpt_pf_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_14_bp_debug_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_14_bp_xcpt_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_14_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_14_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_14_edge_inst = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_14_ftq_idx = 3'b000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_14_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_14_is_rvc = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_14_is_sfb = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_14_pc_lob = 6'b000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_14_taken = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_14_xcpt_ae_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_14_xcpt_pf_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_15_bp_debug_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_15_bp_xcpt_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_15_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_15_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_15_edge_inst = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_15_ftq_idx = 3'b111;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_15_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_15_is_rvc = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_15_is_sfb = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_15_pc_lob = 6'b000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_15_taken = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_15_xcpt_ae_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_15_xcpt_pf_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_1_bp_debug_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_1_bp_xcpt_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_1_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_1_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_1_edge_inst = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_1_ftq_idx = 3'b111;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_1_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_1_is_rvc = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_1_is_sfb = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_1_pc_lob = 6'b000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_1_taken = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_1_xcpt_ae_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_1_xcpt_pf_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_2_bp_debug_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_2_bp_xcpt_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_2_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_2_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_2_edge_inst = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_2_ftq_idx = 3'b000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_2_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_2_is_rvc = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_2_is_sfb = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_2_pc_lob = 6'b000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_2_taken = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_2_xcpt_ae_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_2_xcpt_pf_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_3_bp_debug_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_3_bp_xcpt_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_3_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_3_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_3_edge_inst = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_3_ftq_idx = 3'b111;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_3_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_3_is_rvc = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_3_is_sfb = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_3_pc_lob = 6'b000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_3_taken = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_3_xcpt_ae_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_3_xcpt_pf_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_4_bp_debug_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_4_bp_xcpt_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_4_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_4_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_4_edge_inst = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_4_ftq_idx = 3'b000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_4_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_4_is_rvc = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_4_is_sfb = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_4_pc_lob = 6'b000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_4_taken = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_4_xcpt_ae_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_4_xcpt_pf_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_5_bp_debug_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_5_bp_xcpt_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_5_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_5_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_5_edge_inst = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_5_ftq_idx = 3'b111;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_5_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_5_is_rvc = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_5_is_sfb = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_5_pc_lob = 6'b000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_5_taken = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_5_xcpt_ae_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_5_xcpt_pf_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_6_bp_debug_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_6_bp_xcpt_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_6_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_6_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_6_edge_inst = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_6_ftq_idx = 3'b000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_6_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_6_is_rvc = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_6_is_sfb = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_6_pc_lob = 6'b000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_6_taken = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_6_xcpt_ae_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_6_xcpt_pf_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_7_bp_debug_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_7_bp_xcpt_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_7_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_7_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_7_edge_inst = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_7_ftq_idx = 3'b111;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_7_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_7_is_rvc = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_7_is_sfb = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_7_pc_lob = 6'b000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_7_taken = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_7_xcpt_ae_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_7_xcpt_pf_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_8_bp_debug_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_8_bp_xcpt_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_8_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_8_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_8_edge_inst = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_8_ftq_idx = 3'b000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_8_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_8_is_rvc = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_8_is_sfb = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_8_pc_lob = 6'b000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_8_taken = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_8_xcpt_ae_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_8_xcpt_pf_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_9_bp_debug_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_9_bp_xcpt_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_9_debug_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_9_debug_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_9_edge_inst = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_9_ftq_idx = 3'b111;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_9_inst = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_9_is_rvc = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_9_is_sfb = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_9_pc_lob = 6'b000000;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_9_taken = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_9_xcpt_ae_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.fb_uop_ram_9_xcpt_pf_if = 1'b0;
    UUT.wrapper.uut.frontend.fb.head = 8'b11101111;
    UUT.wrapper.uut.frontend.fb.maybe_full = 1'b0;
    UUT.wrapper.uut.frontend.fb.tail = 16'b0000000001000000;
    UUT.wrapper.uut.frontend.ftq.REG = 1'b0;
    UUT.wrapper.uut.frontend.ftq.REG_1 = 1'b0;
    UUT.wrapper.uut.frontend.ftq.REG_3 = 1'b1;
    UUT.wrapper.uut.frontend.ftq.REG_4 = 3'b111;
    UUT.wrapper.uut.frontend.ftq.bpd_end_idx = 3'b000;
    UUT.wrapper.uut.frontend.ftq.bpd_end_idx_REG = 3'b000;
    UUT.wrapper.uut.frontend.ftq.bpd_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.frontend.ftq.bpd_ptr = 3'b000;
    UUT.wrapper.uut.frontend.ftq.bpd_repair_idx = 3'b000;
    UUT.wrapper.uut.frontend.ftq.bpd_repair_idx_REG = 3'b000;
    UUT.wrapper.uut.frontend.ftq.bpd_repair_pc = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.frontend.ftq.bpd_update_mispredict = 1'b0;
    UUT.wrapper.uut.frontend.ftq.bpd_update_repair = 1'b0;
    UUT.wrapper.uut.frontend.ftq.deq_ptr = 3'b111;
    UUT.wrapper.uut.frontend.ftq.do_commit_update_REG = 1'b0;
    UUT.wrapper.uut.frontend.ftq.enq_ptr = 3'b111;
    UUT.wrapper.uut.frontend.ftq.ghist_0_current_saw_branch_not_taken_bpd_ghist_addr_pipe_0 = 3'b000;
    UUT.wrapper.uut.frontend.ftq.ghist_0_old_history_bpd_ghist_addr_pipe_0 = 3'b000;
    UUT.wrapper.uut.frontend.ftq.ghist_1_current_saw_branch_not_taken_io_get_ftq_pc_1_ghist_MPORT_addr_pipe_0 = 3'b000;
    UUT.wrapper.uut.frontend.ftq.ghist_1_new_saw_branch_not_taken_io_get_ftq_pc_1_ghist_MPORT_addr_pipe_0 = 3'b000;
    UUT.wrapper.uut.frontend.ftq.ghist_1_new_saw_branch_taken_io_get_ftq_pc_1_ghist_MPORT_addr_pipe_0 = 3'b000;
    UUT.wrapper.uut.frontend.ftq.ghist_1_old_history_io_get_ftq_pc_1_ghist_MPORT_addr_pipe_0 = 3'b000;
    UUT.wrapper.uut.frontend.ftq.io_enq_ready_REG = 1'b1;
    UUT.wrapper.uut.frontend.ftq.io_get_ftq_pc_0_com_pc_REG = 40'b0000000000000000000000000000000000111111;
    UUT.wrapper.uut.frontend.ftq.io_get_ftq_pc_0_entry_REG_cfi_idx_bits = 2'b00;
    UUT.wrapper.uut.frontend.ftq.io_get_ftq_pc_0_entry_REG_cfi_idx_valid = 1'b0;
    UUT.wrapper.uut.frontend.ftq.io_get_ftq_pc_0_next_pc_REG = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.frontend.ftq.io_get_ftq_pc_0_next_val_REG = 1'b0;
    UUT.wrapper.uut.frontend.ftq.io_get_ftq_pc_0_pc_REG = 40'b1111111111111111111111111111111011111111;
    UUT.wrapper.uut.frontend.ftq.io_get_ftq_pc_1_entry_REG_br_mask = 4'b0000;
    UUT.wrapper.uut.frontend.ftq.io_get_ftq_pc_1_pc_REG = 40'b0000000000000000000000000000000000111111;
    UUT.wrapper.uut.frontend.ftq.pcs_0 = 40'b0000000000010000000000000000000000000000;
    UUT.wrapper.uut.frontend.ftq.pcs_1 = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.frontend.ftq.pcs_2 = 40'b0000000000000000000000000000000000001000;
    UUT.wrapper.uut.frontend.ftq.pcs_3 = 40'b0000000000010000000000000000000000010000;
    UUT.wrapper.uut.frontend.ftq.pcs_4 = 40'b0000000000010000000000000000000000011000;
    UUT.wrapper.uut.frontend.ftq.pcs_5 = 40'b0000000000010000000000000000000000100000;
    UUT.wrapper.uut.frontend.ftq.pcs_6 = 40'b0000000000010000000000000000000000101000;
    UUT.wrapper.uut.frontend.ftq.pcs_7 = 40'b0000000000000000000000000000000010000000;
    UUT.wrapper.uut.frontend.ftq.prev_entry_REG_br_mask = 4'b0000;
    UUT.wrapper.uut.frontend.ftq.prev_entry_REG_cfi_idx_bits = 2'b00;
    UUT.wrapper.uut.frontend.ftq.prev_entry_REG_cfi_idx_valid = 1'b0;
    UUT.wrapper.uut.frontend.ftq.prev_entry_REG_cfi_taken = 1'b0;
    UUT.wrapper.uut.frontend.ftq.prev_entry_br_mask = 4'b1000;
    UUT.wrapper.uut.frontend.ftq.prev_entry_cfi_idx_bits = 2'b11;
    UUT.wrapper.uut.frontend.ftq.prev_entry_cfi_idx_valid = 1'b1;
    UUT.wrapper.uut.frontend.ftq.prev_entry_cfi_taken = 1'b1;
    UUT.wrapper.uut.frontend.ftq.prev_ghist_current_saw_branch_not_taken = 1'b0;
    UUT.wrapper.uut.frontend.ftq.prev_ghist_old_history = 64'b1110000000000000001111111001100110011001100110011001100110011001;
    UUT.wrapper.uut.frontend.ftq.ram_0_br_mask = 4'b0000;
    UUT.wrapper.uut.frontend.ftq.ram_0_cfi_idx_bits = 2'b11;
    UUT.wrapper.uut.frontend.ftq.ram_0_cfi_idx_valid = 1'b0;
    UUT.wrapper.uut.frontend.ftq.ram_0_cfi_taken = 1'b1;
    UUT.wrapper.uut.frontend.ftq.ram_1_br_mask = 4'b0000;
    UUT.wrapper.uut.frontend.ftq.ram_1_cfi_idx_bits = 2'b00;
    UUT.wrapper.uut.frontend.ftq.ram_1_cfi_idx_valid = 1'b1;
    UUT.wrapper.uut.frontend.ftq.ram_1_cfi_taken = 1'b1;
    UUT.wrapper.uut.frontend.ftq.ram_2_br_mask = 4'b0001;
    UUT.wrapper.uut.frontend.ftq.ram_2_cfi_idx_bits = 2'b00;
    UUT.wrapper.uut.frontend.ftq.ram_2_cfi_idx_valid = 1'b0;
    UUT.wrapper.uut.frontend.ftq.ram_2_cfi_taken = 1'b1;
    UUT.wrapper.uut.frontend.ftq.ram_3_br_mask = 4'b0000;
    UUT.wrapper.uut.frontend.ftq.ram_3_cfi_idx_bits = 2'b11;
    UUT.wrapper.uut.frontend.ftq.ram_3_cfi_idx_valid = 1'b0;
    UUT.wrapper.uut.frontend.ftq.ram_3_cfi_taken = 1'b1;
    UUT.wrapper.uut.frontend.ftq.ram_4_br_mask = 4'b1000;
    UUT.wrapper.uut.frontend.ftq.ram_4_cfi_idx_bits = 2'b11;
    UUT.wrapper.uut.frontend.ftq.ram_4_cfi_idx_valid = 1'b1;
    UUT.wrapper.uut.frontend.ftq.ram_4_cfi_taken = 1'b1;
    UUT.wrapper.uut.frontend.ftq.ram_5_br_mask = 4'b0001;
    UUT.wrapper.uut.frontend.ftq.ram_5_cfi_idx_bits = 2'b11;
    UUT.wrapper.uut.frontend.ftq.ram_5_cfi_idx_valid = 1'b0;
    UUT.wrapper.uut.frontend.ftq.ram_5_cfi_taken = 1'b1;
    UUT.wrapper.uut.frontend.ftq.ram_6_br_mask = 4'b0000;
    UUT.wrapper.uut.frontend.ftq.ram_6_cfi_idx_bits = 2'b11;
    UUT.wrapper.uut.frontend.ftq.ram_6_cfi_idx_valid = 1'b0;
    UUT.wrapper.uut.frontend.ftq.ram_6_cfi_taken = 1'b1;
    UUT.wrapper.uut.frontend.ftq.ram_7_br_mask = 4'b0000;
    UUT.wrapper.uut.frontend.ftq.ram_7_cfi_idx_bits = 2'b00;
    UUT.wrapper.uut.frontend.ftq.ram_7_cfi_idx_valid = 1'b0;
    UUT.wrapper.uut.frontend.ftq.ram_7_cfi_taken = 1'b1;
    UUT.wrapper.uut.frontend.ftq.ram_REG_br_mask = 4'b1111;
    UUT.wrapper.uut.frontend.ftq.ram_REG_cfi_idx_bits = 2'b11;
    UUT.wrapper.uut.frontend.ftq.ram_REG_cfi_idx_valid = 1'b1;
    UUT.wrapper.uut.frontend.ftq.ram_REG_cfi_taken = 1'b1;
    UUT.wrapper.uut.frontend.icache.counter = 3'b001;
    UUT.wrapper.uut.frontend.icache.dataArrayWay_0_s2_dout_0_MPORT_addr_pipe_0 = 4'b1011;
    UUT.wrapper.uut.frontend.icache.invalidated = 1'b0;
    UUT.wrapper.uut.frontend.icache.refill_paddr = 32'b00010000000000000000000011111000;
    UUT.wrapper.uut.frontend.icache.refill_valid = 1'b0;
    UUT.wrapper.uut.frontend.icache.s1_valid = 1'b1;
    UUT.wrapper.uut.frontend.icache.s2_dout_0_REG = 64'b1100001101100001010001110001110110110000011111001111111111111111;
    UUT.wrapper.uut.frontend.icache.s2_hit = 1'b1;
    UUT.wrapper.uut.frontend.icache.s2_miss_REG = 1'b0;
    UUT.wrapper.uut.frontend.icache.s2_valid = 1'b1;
    UUT.wrapper.uut.frontend.icache.tag_array_0_tag_rdata_addr_pipe_0 = 1'b0;
    UUT.wrapper.uut.frontend.icache.vb_array = 2'b11;
    UUT.wrapper.uut.frontend.s1_ghist_current_saw_branch_not_taken = 1'b0;
    UUT.wrapper.uut.frontend.s1_ghist_new_saw_branch_not_taken = 1'b0;
    UUT.wrapper.uut.frontend.s1_ghist_new_saw_branch_taken = 1'b0;
    UUT.wrapper.uut.frontend.s1_ghist_old_history = 64'b1110011001100110011001100110011001100110011001100110011001100101;
    UUT.wrapper.uut.frontend.s1_is_replay = 1'b1;
    UUT.wrapper.uut.frontend.s1_is_sfence = 1'b1;
    UUT.wrapper.uut.frontend.s1_ppc_REG = 32'b00000000000000000000000001111000;
    UUT.wrapper.uut.frontend.s1_tlb_resp_REG_ae_inst = 1'b0;
    UUT.wrapper.uut.frontend.s1_tlb_resp_REG_pf_inst = 1'b0;
    UUT.wrapper.uut.frontend.s1_valid = 1'b1;
    UUT.wrapper.uut.frontend.s1_vpc = 40'b0011111111011101111000000000000000000000;
    UUT.wrapper.uut.frontend.s2_ghist_current_saw_branch_not_taken = 1'b1;
    UUT.wrapper.uut.frontend.s2_ghist_new_saw_branch_not_taken = 1'b0;
    UUT.wrapper.uut.frontend.s2_ghist_new_saw_branch_taken = 1'b0;
    UUT.wrapper.uut.frontend.s2_ghist_old_history = 64'b1110011001100110011001100110011001100110011001100110011001100101;
    UUT.wrapper.uut.frontend.s2_is_replay_REG = 1'b1;
    UUT.wrapper.uut.frontend.s2_ppc = 32'b00010000000000000000100000111000;
    UUT.wrapper.uut.frontend.s2_tlb_miss = 1'b0;
    UUT.wrapper.uut.frontend.s2_tlb_resp_ae_inst = 1'b1;
    UUT.wrapper.uut.frontend.s2_tlb_resp_pf_inst = 1'b1;
    UUT.wrapper.uut.frontend.s2_valid = 1'b1;
    UUT.wrapper.uut.frontend.s2_vpc = 40'b0011111111011101111000000000000000000000;
    UUT.wrapper.uut.frontend.tlb.r_need_gpa = 1'b0;
    UUT.wrapper.uut.frontend.tlb.r_refill_tag = 27'b000000000010000000000000000;
    UUT.wrapper.uut.frontend.tlb.r_sectored_hit_valid = 1'b1;
    UUT.wrapper.uut.frontend.tlb.r_superpage_repl_addr = 2'b11;
    UUT.wrapper.uut.frontend.tlb.sectored_entries_0_0_data_0 = 42'b000000000000000000000010001000111101111111;
    UUT.wrapper.uut.frontend.tlb.sectored_entries_0_0_data_1 = 42'b000000000000000000000000001000111101111111;
    UUT.wrapper.uut.frontend.tlb.sectored_entries_0_0_data_2 = 42'b000000000000000000000000101101111101111111;
    UUT.wrapper.uut.frontend.tlb.sectored_entries_0_0_data_3 = 42'b000000000000000000000000001000111001000011;
    UUT.wrapper.uut.frontend.tlb.sectored_entries_0_0_tag_vpn = 27'b000000000000000000000000000;
    UUT.wrapper.uut.frontend.tlb.sectored_entries_0_0_valid_0 = 1'b0;
    UUT.wrapper.uut.frontend.tlb.sectored_entries_0_0_valid_1 = 1'b1;
    UUT.wrapper.uut.frontend.tlb.sectored_entries_0_0_valid_2 = 1'b1;
    UUT.wrapper.uut.frontend.tlb.sectored_entries_0_0_valid_3 = 1'b0;
    UUT.wrapper.uut.frontend.tlb.special_entry_data_0 = 42'b000000000000000011110010011000111100100001;
    UUT.wrapper.uut.frontend.tlb.special_entry_level = 2'b10;
    UUT.wrapper.uut.frontend.tlb.special_entry_tag_vpn = 27'b011111111011101111000000000;
    UUT.wrapper.uut.frontend.tlb.special_entry_valid_0 = 1'b1;
    UUT.wrapper.uut.frontend.tlb.state = 2'b01;
    UUT.wrapper.uut.frontend.tlb.state_reg_1 = 3'b010;
    UUT.wrapper.uut.frontend.tlb.superpage_entries_0_data_0 = 42'b000000000000000000000010001101111101111111;
    UUT.wrapper.uut.frontend.tlb.superpage_entries_0_level = 2'b00;
    UUT.wrapper.uut.frontend.tlb.superpage_entries_0_tag_vpn = 27'b000000000010000000000000011;
    UUT.wrapper.uut.frontend.tlb.superpage_entries_0_valid_0 = 1'b1;
    UUT.wrapper.uut.frontend.tlb.superpage_entries_1_data_0 = 42'b000000000000000000000010101101111101111111;
    UUT.wrapper.uut.frontend.tlb.superpage_entries_1_level = 2'b00;
    UUT.wrapper.uut.frontend.tlb.superpage_entries_1_tag_vpn = 27'b000000000010000000000000000;
    UUT.wrapper.uut.frontend.tlb.superpage_entries_1_valid_0 = 1'b1;
    UUT.wrapper.uut.frontend.tlb.superpage_entries_2_data_0 = 42'b000000000000000000000010101101111101111111;
    UUT.wrapper.uut.frontend.tlb.superpage_entries_2_level = 2'b00;
    UUT.wrapper.uut.frontend.tlb.superpage_entries_2_tag_vpn = 27'b000000000010000000000000000;
    UUT.wrapper.uut.frontend.tlb.superpage_entries_2_valid_0 = 1'b1;
    UUT.wrapper.uut.frontend.tlb.superpage_entries_3_data_0 = 42'b000000000000000000000010101101111101111111;
    UUT.wrapper.uut.frontend.tlb.superpage_entries_3_level = 2'b00;
    UUT.wrapper.uut.frontend.tlb.superpage_entries_3_tag_vpn = 27'b000000000010000000000000000;
    UUT.wrapper.uut.frontend.tlb.superpage_entries_3_valid_0 = 1'b1;
    UUT.wrapper.uut.frontend.tlb_io_sfence_REG_bits_addr = 39'b000000000000000000000000000000000000000;
    UUT.wrapper.uut.frontend.tlb_io_sfence_REG_bits_rs1 = 1'b0;
    UUT.wrapper.uut.frontend.tlb_io_sfence_REG_bits_rs2 = 1'b0;
    UUT.wrapper.uut.frontend.tlb_io_sfence_REG_valid = 1'b0;
    UUT.wrapper.uut.lsu.REG = 1'b0;
    UUT.wrapper.uut.lsu.REG_1 = 1'b0;
    UUT.wrapper.uut.lsu.can_fire_load_retry_REG = 1'b1;
    UUT.wrapper.uut.lsu.can_fire_sta_retry_REG = 1'b0;
    UUT.wrapper.uut.lsu.clr_bsy_brmask_0 = 12'b000000000000;
    UUT.wrapper.uut.lsu.clr_bsy_rob_idx_0 = 6'b000000;
    UUT.wrapper.uut.lsu.clr_bsy_valid_0 = 1'b0;
    UUT.wrapper.uut.lsu.dtlb.r_refill_tag = 27'b111111111111111111111111111;
    UUT.wrapper.uut.lsu.dtlb.r_sectored_hit = 1'b0;
    UUT.wrapper.uut.lsu.dtlb.r_superpage_repl_addr = 2'b11;
    UUT.wrapper.uut.lsu.dtlb.sectored_entries_0_data_0 = 34'b0000000000000000000000000001000001;
    UUT.wrapper.uut.lsu.dtlb.sectored_entries_0_data_1 = 34'b0000000000000000000011111111111111;
    UUT.wrapper.uut.lsu.dtlb.sectored_entries_0_data_2 = 34'b1111111111100000000010101111111110;
    UUT.wrapper.uut.lsu.dtlb.sectored_entries_0_data_3 = 34'b0000001000000000000011111110111110;
    UUT.wrapper.uut.lsu.dtlb.sectored_entries_0_tag = 27'b011111111111111111111111100;
    UUT.wrapper.uut.lsu.dtlb.sectored_entries_0_valid_0 = 1'b1;
    UUT.wrapper.uut.lsu.dtlb.sectored_entries_0_valid_1 = 1'b1;
    UUT.wrapper.uut.lsu.dtlb.sectored_entries_0_valid_2 = 1'b1;
    UUT.wrapper.uut.lsu.dtlb.sectored_entries_0_valid_3 = 1'b1;
    UUT.wrapper.uut.lsu.dtlb.special_entry_data_0 = 34'b0000000000000000000010100011100010;
    UUT.wrapper.uut.lsu.dtlb.special_entry_level = 2'b00;
    UUT.wrapper.uut.lsu.dtlb.special_entry_tag = 27'b001100111000000000000000000;
    UUT.wrapper.uut.lsu.dtlb.special_entry_valid_0 = 1'b1;
    UUT.wrapper.uut.lsu.dtlb.state = 2'b01;
    UUT.wrapper.uut.lsu.dtlb.state_reg_1 = 3'b000;
    UUT.wrapper.uut.lsu.dtlb.superpage_entries_0_data_0 = 34'b0000000000000000000000000001000001;
    UUT.wrapper.uut.lsu.dtlb.superpage_entries_0_level = 2'b00;
    UUT.wrapper.uut.lsu.dtlb.superpage_entries_0_tag = 27'b011111111000000000111111111;
    UUT.wrapper.uut.lsu.dtlb.superpage_entries_0_valid_0 = 1'b1;
    UUT.wrapper.uut.lsu.dtlb.superpage_entries_1_data_0 = 34'b1111111111111111111101011111111001;
    UUT.wrapper.uut.lsu.dtlb.superpage_entries_1_level = 2'b10;
    UUT.wrapper.uut.lsu.dtlb.superpage_entries_1_tag = 27'b001100111111111111111111111;
    UUT.wrapper.uut.lsu.dtlb.superpage_entries_1_valid_0 = 1'b1;
    UUT.wrapper.uut.lsu.dtlb.superpage_entries_2_data_0 = 34'b0000000000011111111101010111111001;
    UUT.wrapper.uut.lsu.dtlb.superpage_entries_2_level = 2'b10;
    UUT.wrapper.uut.lsu.dtlb.superpage_entries_2_tag = 27'b001100111111111111111111111;
    UUT.wrapper.uut.lsu.dtlb.superpage_entries_2_valid_0 = 1'b1;
    UUT.wrapper.uut.lsu.dtlb.superpage_entries_3_data_0 = 34'b0000000000011111111101010111111001;
    UUT.wrapper.uut.lsu.dtlb.superpage_entries_3_level = 2'b10;
    UUT.wrapper.uut.lsu.dtlb.superpage_entries_3_tag = 27'b001100111111111111111111111;
    UUT.wrapper.uut.lsu.dtlb.superpage_entries_3_valid_0 = 1'b1;
    UUT.wrapper.uut.lsu.fired_load_incoming_REG = 1'b1;
    UUT.wrapper.uut.lsu.fired_load_retry_REG = 1'b0;
    UUT.wrapper.uut.lsu.fired_load_wakeup_REG = 1'b0;
    UUT.wrapper.uut.lsu.fired_release_0 = 1'b1;
    UUT.wrapper.uut.lsu.fired_sfence_0 = 1'b0;
    UUT.wrapper.uut.lsu.fired_sta_incoming_REG = 1'b0;
    UUT.wrapper.uut.lsu.fired_sta_retry_REG = 1'b0;
    UUT.wrapper.uut.lsu.fired_stad_incoming_REG = 1'b0;
    UUT.wrapper.uut.lsu.fired_std_incoming_REG = 1'b0;
    UUT.wrapper.uut.lsu.hella_paddr = 32'b00000000000000000000000000000000;
    UUT.wrapper.uut.lsu.hella_req_addr = 40'b1111111100000000000000000000000001111000;
    UUT.wrapper.uut.lsu.hella_state = 3'b100;
    UUT.wrapper.uut.lsu.hella_xcpt_ae_ld = 1'b1;
    UUT.wrapper.uut.lsu.hella_xcpt_ae_st = 1'b0;
    UUT.wrapper.uut.lsu.hella_xcpt_ma_ld = 1'b0;
    UUT.wrapper.uut.lsu.hella_xcpt_ma_st = 1'b0;
    UUT.wrapper.uut.lsu.hella_xcpt_pf_ld = 1'b0;
    UUT.wrapper.uut.lsu.hella_xcpt_pf_st = 1'b0;
    UUT.wrapper.uut.lsu.io_core_clr_bsy_0_valid_REG = 1'b0;
    UUT.wrapper.uut.lsu.io_core_clr_bsy_0_valid_REG_1 = 1'b0;
    UUT.wrapper.uut.lsu.io_core_clr_bsy_0_valid_REG_2 = 1'b0;
    UUT.wrapper.uut.lsu.io_core_ld_miss_REG = 1'b1;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG = 1'b0;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_1 = 1'b1;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_10 = 1'b1;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_11 = 1'b0;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_12 = 1'b0;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_13 = 1'b0;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_14 = 1'b0;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_15 = 1'b1;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_16 = 1'b0;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_17 = 1'b0;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_18 = 1'b0;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_19 = 1'b1;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_2 = 1'b1;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_20 = 1'b1;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_21 = 1'b1;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_22 = 1'b0;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_23 = 1'b0;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_24 = 1'b0;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_25 = 1'b1;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_26 = 1'b1;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_27 = 1'b1;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_28 = 1'b1;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_29 = 1'b0;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_3 = 1'b1;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_30 = 1'b0;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_31 = 1'b1;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_32 = 1'b1;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_33 = 1'b1;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_34 = 1'b1;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_35 = 1'b1;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_36 = 1'b0;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_37 = 1'b1;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_38 = 1'b1;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_39 = 1'b1;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_4 = 1'b1;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_40 = 1'b0;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_41 = 1'b1;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_42 = 1'b0;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_43 = 1'b1;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_44 = 1'b1;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_45 = 1'b1;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_46 = 1'b0;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_47 = 1'b0;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_48 = 1'b0;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_49 = 1'b1;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_5 = 1'b1;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_50 = 1'b1;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_51 = 1'b1;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_52 = 1'b0;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_53 = 1'b1;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_54 = 1'b0;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_55 = 1'b1;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_56 = 1'b1;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_57 = 1'b1;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_58 = 1'b0;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_59 = 1'b1;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_6 = 1'b1;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_60 = 1'b1;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_61 = 1'b0;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_62 = 1'b0;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_63 = 1'b0;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_7 = 1'b1;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_8 = 1'b1;
    UUT.wrapper.uut.lsu.io_dmem_s1_kill_0_REG_9 = 1'b1;
    UUT.wrapper.uut.lsu.lcam_addr_REG = 32'b00000000000000000000000000000100;
    UUT.wrapper.uut.lsu.lcam_addr_REG_1 = 32'b10000000000000000000000000000110;
    UUT.wrapper.uut.lsu.lcam_ldq_idx_REG = 4'b0000;
    UUT.wrapper.uut.lsu.lcam_ldq_idx_REG_1 = 4'b1111;
    UUT.wrapper.uut.lsu.lcam_stq_idx_REG = 4'b1010;
    UUT.wrapper.uut.lsu.ldq_0_bits_addr_bits = 40'b0000000000011101100110011001100000010001;
    UUT.wrapper.uut.lsu.ldq_0_bits_addr_is_uncacheable = 1'b0;
    UUT.wrapper.uut.lsu.ldq_0_bits_addr_is_virtual = 1'b0;
    UUT.wrapper.uut.lsu.ldq_0_bits_addr_valid = 1'b1;
    UUT.wrapper.uut.lsu.ldq_0_bits_debug_wb_data = 64'b0000000000000000000000000000000000000000000000000000000010100000;
    UUT.wrapper.uut.lsu.ldq_0_bits_executed = 1'b1;
    UUT.wrapper.uut.lsu.ldq_0_bits_forward_std_val = 1'b0;
    UUT.wrapper.uut.lsu.ldq_0_bits_forward_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_0_bits_observed = 1'b0;
    UUT.wrapper.uut.lsu.ldq_0_bits_order_fail = 1'b1;
    UUT.wrapper.uut.lsu.ldq_0_bits_st_dep_mask = 16'b0000000000000000;
    UUT.wrapper.uut.lsu.ldq_0_bits_succeeded = 1'b0;
    UUT.wrapper.uut.lsu.ldq_0_bits_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.lsu.ldq_0_bits_uop_dst_rtype = 2'b00;
    UUT.wrapper.uut.lsu.ldq_0_bits_uop_is_amo = 1'b0;
    UUT.wrapper.uut.lsu.ldq_0_bits_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_0_bits_uop_mem_cmd = 5'b00000;
    UUT.wrapper.uut.lsu.ldq_0_bits_uop_mem_signed = 1'b0;
    UUT.wrapper.uut.lsu.ldq_0_bits_uop_mem_size = 2'b11;
    UUT.wrapper.uut.lsu.ldq_0_bits_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.lsu.ldq_0_bits_uop_rob_idx = 6'b000011;
    UUT.wrapper.uut.lsu.ldq_0_bits_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_0_bits_uop_uses_ldq = 1'b1;
    UUT.wrapper.uut.lsu.ldq_0_bits_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.lsu.ldq_0_bits_youngest_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_0_valid = 1'b1;
    UUT.wrapper.uut.lsu.ldq_10_bits_addr_bits = 40'b0001100111111111111111111111100111011111;
    UUT.wrapper.uut.lsu.ldq_10_bits_addr_is_uncacheable = 1'b1;
    UUT.wrapper.uut.lsu.ldq_10_bits_addr_is_virtual = 1'b1;
    UUT.wrapper.uut.lsu.ldq_10_bits_addr_valid = 1'b1;
    UUT.wrapper.uut.lsu.ldq_10_bits_debug_wb_data = 64'b1111111111111111111111111111111111111111111111111111111111111111;
    UUT.wrapper.uut.lsu.ldq_10_bits_executed = 1'b1;
    UUT.wrapper.uut.lsu.ldq_10_bits_forward_std_val = 1'b1;
    UUT.wrapper.uut.lsu.ldq_10_bits_forward_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_10_bits_observed = 1'b0;
    UUT.wrapper.uut.lsu.ldq_10_bits_order_fail = 1'b1;
    UUT.wrapper.uut.lsu.ldq_10_bits_st_dep_mask = 16'b1111111111111110;
    UUT.wrapper.uut.lsu.ldq_10_bits_succeeded = 1'b1;
    UUT.wrapper.uut.lsu.ldq_10_bits_uop_br_mask = 12'b111100000000;
    UUT.wrapper.uut.lsu.ldq_10_bits_uop_dst_rtype = 2'b11;
    UUT.wrapper.uut.lsu.ldq_10_bits_uop_is_amo = 1'b1;
    UUT.wrapper.uut.lsu.ldq_10_bits_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_10_bits_uop_mem_cmd = 5'b00000;
    UUT.wrapper.uut.lsu.ldq_10_bits_uop_mem_signed = 1'b1;
    UUT.wrapper.uut.lsu.ldq_10_bits_uop_mem_size = 2'b11;
    UUT.wrapper.uut.lsu.ldq_10_bits_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.lsu.ldq_10_bits_uop_rob_idx = 6'b000000;
    UUT.wrapper.uut.lsu.ldq_10_bits_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_10_bits_uop_uses_ldq = 1'b1;
    UUT.wrapper.uut.lsu.ldq_10_bits_uop_uses_stq = 1'b1;
    UUT.wrapper.uut.lsu.ldq_10_bits_youngest_stq_idx = 4'b1111;
    UUT.wrapper.uut.lsu.ldq_10_valid = 1'b0;
    UUT.wrapper.uut.lsu.ldq_11_bits_addr_bits = 40'b0001100111111111111111111111100111011111;
    UUT.wrapper.uut.lsu.ldq_11_bits_addr_is_uncacheable = 1'b1;
    UUT.wrapper.uut.lsu.ldq_11_bits_addr_is_virtual = 1'b1;
    UUT.wrapper.uut.lsu.ldq_11_bits_addr_valid = 1'b1;
    UUT.wrapper.uut.lsu.ldq_11_bits_debug_wb_data = 64'b1111111111111111111111111111111111111111111111111111111111111111;
    UUT.wrapper.uut.lsu.ldq_11_bits_executed = 1'b1;
    UUT.wrapper.uut.lsu.ldq_11_bits_forward_std_val = 1'b1;
    UUT.wrapper.uut.lsu.ldq_11_bits_forward_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_11_bits_observed = 1'b0;
    UUT.wrapper.uut.lsu.ldq_11_bits_order_fail = 1'b1;
    UUT.wrapper.uut.lsu.ldq_11_bits_st_dep_mask = 16'b1111111111111110;
    UUT.wrapper.uut.lsu.ldq_11_bits_succeeded = 1'b1;
    UUT.wrapper.uut.lsu.ldq_11_bits_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.lsu.ldq_11_bits_uop_dst_rtype = 2'b11;
    UUT.wrapper.uut.lsu.ldq_11_bits_uop_is_amo = 1'b1;
    UUT.wrapper.uut.lsu.ldq_11_bits_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_11_bits_uop_mem_cmd = 5'b00000;
    UUT.wrapper.uut.lsu.ldq_11_bits_uop_mem_signed = 1'b1;
    UUT.wrapper.uut.lsu.ldq_11_bits_uop_mem_size = 2'b11;
    UUT.wrapper.uut.lsu.ldq_11_bits_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.lsu.ldq_11_bits_uop_rob_idx = 6'b000000;
    UUT.wrapper.uut.lsu.ldq_11_bits_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_11_bits_uop_uses_ldq = 1'b1;
    UUT.wrapper.uut.lsu.ldq_11_bits_uop_uses_stq = 1'b1;
    UUT.wrapper.uut.lsu.ldq_11_bits_youngest_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_11_valid = 1'b1;
    UUT.wrapper.uut.lsu.ldq_12_bits_addr_bits = 40'b0001100110011001100110011001100111011110;
    UUT.wrapper.uut.lsu.ldq_12_bits_addr_is_uncacheable = 1'b1;
    UUT.wrapper.uut.lsu.ldq_12_bits_addr_is_virtual = 1'b1;
    UUT.wrapper.uut.lsu.ldq_12_bits_addr_valid = 1'b1;
    UUT.wrapper.uut.lsu.ldq_12_bits_debug_wb_data = 64'b0000000000000000000000000000000000000000000000001000000010000000;
    UUT.wrapper.uut.lsu.ldq_12_bits_executed = 1'b1;
    UUT.wrapper.uut.lsu.ldq_12_bits_forward_std_val = 1'b1;
    UUT.wrapper.uut.lsu.ldq_12_bits_forward_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_12_bits_observed = 1'b0;
    UUT.wrapper.uut.lsu.ldq_12_bits_order_fail = 1'b1;
    UUT.wrapper.uut.lsu.ldq_12_bits_st_dep_mask = 16'b1111111111111110;
    UUT.wrapper.uut.lsu.ldq_12_bits_succeeded = 1'b1;
    UUT.wrapper.uut.lsu.ldq_12_bits_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.lsu.ldq_12_bits_uop_dst_rtype = 2'b11;
    UUT.wrapper.uut.lsu.ldq_12_bits_uop_is_amo = 1'b1;
    UUT.wrapper.uut.lsu.ldq_12_bits_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_12_bits_uop_mem_cmd = 5'b00000;
    UUT.wrapper.uut.lsu.ldq_12_bits_uop_mem_signed = 1'b1;
    UUT.wrapper.uut.lsu.ldq_12_bits_uop_mem_size = 2'b11;
    UUT.wrapper.uut.lsu.ldq_12_bits_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.lsu.ldq_12_bits_uop_rob_idx = 6'b000000;
    UUT.wrapper.uut.lsu.ldq_12_bits_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_12_bits_uop_uses_ldq = 1'b1;
    UUT.wrapper.uut.lsu.ldq_12_bits_uop_uses_stq = 1'b1;
    UUT.wrapper.uut.lsu.ldq_12_bits_youngest_stq_idx = 4'b1111;
    UUT.wrapper.uut.lsu.ldq_12_valid = 1'b1;
    UUT.wrapper.uut.lsu.ldq_13_bits_addr_bits = 40'b0001100111111111111111111111100111011111;
    UUT.wrapper.uut.lsu.ldq_13_bits_addr_is_uncacheable = 1'b1;
    UUT.wrapper.uut.lsu.ldq_13_bits_addr_is_virtual = 1'b1;
    UUT.wrapper.uut.lsu.ldq_13_bits_addr_valid = 1'b1;
    UUT.wrapper.uut.lsu.ldq_13_bits_debug_wb_data = 64'b1111111111111111111111111111111111111111111111111111111111111111;
    UUT.wrapper.uut.lsu.ldq_13_bits_executed = 1'b1;
    UUT.wrapper.uut.lsu.ldq_13_bits_forward_std_val = 1'b1;
    UUT.wrapper.uut.lsu.ldq_13_bits_forward_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_13_bits_observed = 1'b0;
    UUT.wrapper.uut.lsu.ldq_13_bits_order_fail = 1'b1;
    UUT.wrapper.uut.lsu.ldq_13_bits_st_dep_mask = 16'b1111111111111010;
    UUT.wrapper.uut.lsu.ldq_13_bits_succeeded = 1'b1;
    UUT.wrapper.uut.lsu.ldq_13_bits_uop_br_mask = 12'b110000000000;
    UUT.wrapper.uut.lsu.ldq_13_bits_uop_dst_rtype = 2'b11;
    UUT.wrapper.uut.lsu.ldq_13_bits_uop_is_amo = 1'b1;
    UUT.wrapper.uut.lsu.ldq_13_bits_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_13_bits_uop_mem_cmd = 5'b00000;
    UUT.wrapper.uut.lsu.ldq_13_bits_uop_mem_signed = 1'b1;
    UUT.wrapper.uut.lsu.ldq_13_bits_uop_mem_size = 2'b11;
    UUT.wrapper.uut.lsu.ldq_13_bits_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.lsu.ldq_13_bits_uop_rob_idx = 6'b000000;
    UUT.wrapper.uut.lsu.ldq_13_bits_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_13_bits_uop_uses_ldq = 1'b1;
    UUT.wrapper.uut.lsu.ldq_13_bits_uop_uses_stq = 1'b1;
    UUT.wrapper.uut.lsu.ldq_13_bits_youngest_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_13_valid = 1'b1;
    UUT.wrapper.uut.lsu.ldq_14_bits_addr_bits = 40'b0000100111111111111111111111100111011000;
    UUT.wrapper.uut.lsu.ldq_14_bits_addr_is_uncacheable = 1'b1;
    UUT.wrapper.uut.lsu.ldq_14_bits_addr_is_virtual = 1'b1;
    UUT.wrapper.uut.lsu.ldq_14_bits_addr_valid = 1'b1;
    UUT.wrapper.uut.lsu.ldq_14_bits_debug_wb_data = 64'b1111111111111111111111111111111111111111111111111111111111111111;
    UUT.wrapper.uut.lsu.ldq_14_bits_executed = 1'b1;
    UUT.wrapper.uut.lsu.ldq_14_bits_forward_std_val = 1'b1;
    UUT.wrapper.uut.lsu.ldq_14_bits_forward_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_14_bits_observed = 1'b0;
    UUT.wrapper.uut.lsu.ldq_14_bits_order_fail = 1'b1;
    UUT.wrapper.uut.lsu.ldq_14_bits_st_dep_mask = 16'b1111111111111110;
    UUT.wrapper.uut.lsu.ldq_14_bits_succeeded = 1'b1;
    UUT.wrapper.uut.lsu.ldq_14_bits_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.lsu.ldq_14_bits_uop_dst_rtype = 2'b11;
    UUT.wrapper.uut.lsu.ldq_14_bits_uop_is_amo = 1'b1;
    UUT.wrapper.uut.lsu.ldq_14_bits_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_14_bits_uop_mem_cmd = 5'b00000;
    UUT.wrapper.uut.lsu.ldq_14_bits_uop_mem_signed = 1'b1;
    UUT.wrapper.uut.lsu.ldq_14_bits_uop_mem_size = 2'b00;
    UUT.wrapper.uut.lsu.ldq_14_bits_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.lsu.ldq_14_bits_uop_rob_idx = 6'b000000;
    UUT.wrapper.uut.lsu.ldq_14_bits_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_14_bits_uop_uses_ldq = 1'b1;
    UUT.wrapper.uut.lsu.ldq_14_bits_uop_uses_stq = 1'b1;
    UUT.wrapper.uut.lsu.ldq_14_bits_youngest_stq_idx = 4'b1111;
    UUT.wrapper.uut.lsu.ldq_14_valid = 1'b1;
    UUT.wrapper.uut.lsu.ldq_15_bits_addr_bits = 40'b0001100111111111111111111111100111011111;
    UUT.wrapper.uut.lsu.ldq_15_bits_addr_is_uncacheable = 1'b1;
    UUT.wrapper.uut.lsu.ldq_15_bits_addr_is_virtual = 1'b1;
    UUT.wrapper.uut.lsu.ldq_15_bits_addr_valid = 1'b1;
    UUT.wrapper.uut.lsu.ldq_15_bits_debug_wb_data = 64'b1111111111111111111111111111111111111111111111111111111111111111;
    UUT.wrapper.uut.lsu.ldq_15_bits_executed = 1'b0;
    UUT.wrapper.uut.lsu.ldq_15_bits_forward_std_val = 1'b0;
    UUT.wrapper.uut.lsu.ldq_15_bits_forward_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_15_bits_observed = 1'b0;
    UUT.wrapper.uut.lsu.ldq_15_bits_order_fail = 1'b0;
    UUT.wrapper.uut.lsu.ldq_15_bits_st_dep_mask = 16'b0000000000000000;
    UUT.wrapper.uut.lsu.ldq_15_bits_succeeded = 1'b0;
    UUT.wrapper.uut.lsu.ldq_15_bits_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.lsu.ldq_15_bits_uop_dst_rtype = 2'b11;
    UUT.wrapper.uut.lsu.ldq_15_bits_uop_is_amo = 1'b1;
    UUT.wrapper.uut.lsu.ldq_15_bits_uop_ldq_idx = 4'b1111;
    UUT.wrapper.uut.lsu.ldq_15_bits_uop_mem_cmd = 5'b11111;
    UUT.wrapper.uut.lsu.ldq_15_bits_uop_mem_signed = 1'b1;
    UUT.wrapper.uut.lsu.ldq_15_bits_uop_mem_size = 2'b11;
    UUT.wrapper.uut.lsu.ldq_15_bits_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.lsu.ldq_15_bits_uop_rob_idx = 6'b111111;
    UUT.wrapper.uut.lsu.ldq_15_bits_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_15_bits_uop_uses_ldq = 1'b1;
    UUT.wrapper.uut.lsu.ldq_15_bits_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.lsu.ldq_15_bits_youngest_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_15_valid = 1'b1;
    UUT.wrapper.uut.lsu.ldq_1_bits_addr_bits = 40'b0000000101100110011001100110000111011011;
    UUT.wrapper.uut.lsu.ldq_1_bits_addr_is_uncacheable = 1'b1;
    UUT.wrapper.uut.lsu.ldq_1_bits_addr_is_virtual = 1'b0;
    UUT.wrapper.uut.lsu.ldq_1_bits_addr_valid = 1'b1;
    UUT.wrapper.uut.lsu.ldq_1_bits_debug_wb_data = 64'b0000000000000000000000000000000000000000000000001000000010000000;
    UUT.wrapper.uut.lsu.ldq_1_bits_executed = 1'b1;
    UUT.wrapper.uut.lsu.ldq_1_bits_forward_std_val = 1'b0;
    UUT.wrapper.uut.lsu.ldq_1_bits_forward_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_1_bits_observed = 1'b0;
    UUT.wrapper.uut.lsu.ldq_1_bits_order_fail = 1'b0;
    UUT.wrapper.uut.lsu.ldq_1_bits_st_dep_mask = 16'b0000000000000000;
    UUT.wrapper.uut.lsu.ldq_1_bits_succeeded = 1'b0;
    UUT.wrapper.uut.lsu.ldq_1_bits_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.lsu.ldq_1_bits_uop_dst_rtype = 2'b00;
    UUT.wrapper.uut.lsu.ldq_1_bits_uop_is_amo = 1'b0;
    UUT.wrapper.uut.lsu.ldq_1_bits_uop_ldq_idx = 4'b0001;
    UUT.wrapper.uut.lsu.ldq_1_bits_uop_mem_cmd = 5'b00000;
    UUT.wrapper.uut.lsu.ldq_1_bits_uop_mem_signed = 1'b0;
    UUT.wrapper.uut.lsu.ldq_1_bits_uop_mem_size = 2'b10;
    UUT.wrapper.uut.lsu.ldq_1_bits_uop_pdst = 7'b0000100;
    UUT.wrapper.uut.lsu.ldq_1_bits_uop_rob_idx = 6'b000110;
    UUT.wrapper.uut.lsu.ldq_1_bits_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_1_bits_uop_uses_ldq = 1'b1;
    UUT.wrapper.uut.lsu.ldq_1_bits_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.lsu.ldq_1_bits_youngest_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_1_valid = 1'b1;
    UUT.wrapper.uut.lsu.ldq_2_bits_addr_bits = 40'b0000000001111111111111111111100111011111;
    UUT.wrapper.uut.lsu.ldq_2_bits_addr_is_uncacheable = 1'b1;
    UUT.wrapper.uut.lsu.ldq_2_bits_addr_is_virtual = 1'b0;
    UUT.wrapper.uut.lsu.ldq_2_bits_addr_valid = 1'b1;
    UUT.wrapper.uut.lsu.ldq_2_bits_debug_wb_data = 64'b1111111111111111111111111111111111111111111111111111111111111111;
    UUT.wrapper.uut.lsu.ldq_2_bits_executed = 1'b1;
    UUT.wrapper.uut.lsu.ldq_2_bits_forward_std_val = 1'b0;
    UUT.wrapper.uut.lsu.ldq_2_bits_forward_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_2_bits_observed = 1'b1;
    UUT.wrapper.uut.lsu.ldq_2_bits_order_fail = 1'b0;
    UUT.wrapper.uut.lsu.ldq_2_bits_st_dep_mask = 16'b0000000000000011;
    UUT.wrapper.uut.lsu.ldq_2_bits_succeeded = 1'b0;
    UUT.wrapper.uut.lsu.ldq_2_bits_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.lsu.ldq_2_bits_uop_dst_rtype = 2'b00;
    UUT.wrapper.uut.lsu.ldq_2_bits_uop_is_amo = 1'b0;
    UUT.wrapper.uut.lsu.ldq_2_bits_uop_ldq_idx = 4'b0010;
    UUT.wrapper.uut.lsu.ldq_2_bits_uop_mem_cmd = 5'b00000;
    UUT.wrapper.uut.lsu.ldq_2_bits_uop_mem_signed = 1'b1;
    UUT.wrapper.uut.lsu.ldq_2_bits_uop_mem_size = 2'b11;
    UUT.wrapper.uut.lsu.ldq_2_bits_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.lsu.ldq_2_bits_uop_rob_idx = 6'b000010;
    UUT.wrapper.uut.lsu.ldq_2_bits_uop_stq_idx = 4'b0010;
    UUT.wrapper.uut.lsu.ldq_2_bits_uop_uses_ldq = 1'b1;
    UUT.wrapper.uut.lsu.ldq_2_bits_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.lsu.ldq_2_bits_youngest_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_2_valid = 1'b1;
    UUT.wrapper.uut.lsu.ldq_3_bits_addr_bits = 40'b0000000000000000000000000000000111011011;
    UUT.wrapper.uut.lsu.ldq_3_bits_addr_is_uncacheable = 1'b0;
    UUT.wrapper.uut.lsu.ldq_3_bits_addr_is_virtual = 1'b1;
    UUT.wrapper.uut.lsu.ldq_3_bits_addr_valid = 1'b1;
    UUT.wrapper.uut.lsu.ldq_3_bits_debug_wb_data = 64'b1111111111111111111111111111111111111111111111111111111110000000;
    UUT.wrapper.uut.lsu.ldq_3_bits_executed = 1'b1;
    UUT.wrapper.uut.lsu.ldq_3_bits_forward_std_val = 1'b0;
    UUT.wrapper.uut.lsu.ldq_3_bits_forward_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_3_bits_observed = 1'b1;
    UUT.wrapper.uut.lsu.ldq_3_bits_order_fail = 1'b1;
    UUT.wrapper.uut.lsu.ldq_3_bits_st_dep_mask = 16'b0000000000000001;
    UUT.wrapper.uut.lsu.ldq_3_bits_succeeded = 1'b0;
    UUT.wrapper.uut.lsu.ldq_3_bits_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.lsu.ldq_3_bits_uop_dst_rtype = 2'b01;
    UUT.wrapper.uut.lsu.ldq_3_bits_uop_is_amo = 1'b0;
    UUT.wrapper.uut.lsu.ldq_3_bits_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_3_bits_uop_mem_cmd = 5'b00000;
    UUT.wrapper.uut.lsu.ldq_3_bits_uop_mem_signed = 1'b0;
    UUT.wrapper.uut.lsu.ldq_3_bits_uop_mem_size = 2'b10;
    UUT.wrapper.uut.lsu.ldq_3_bits_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.lsu.ldq_3_bits_uop_rob_idx = 6'b001000;
    UUT.wrapper.uut.lsu.ldq_3_bits_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_3_bits_uop_uses_ldq = 1'b1;
    UUT.wrapper.uut.lsu.ldq_3_bits_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.lsu.ldq_3_bits_youngest_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_3_valid = 1'b1;
    UUT.wrapper.uut.lsu.ldq_4_bits_addr_bits = 40'b0001100111111111111111111111100111011111;
    UUT.wrapper.uut.lsu.ldq_4_bits_addr_is_uncacheable = 1'b1;
    UUT.wrapper.uut.lsu.ldq_4_bits_addr_is_virtual = 1'b1;
    UUT.wrapper.uut.lsu.ldq_4_bits_addr_valid = 1'b1;
    UUT.wrapper.uut.lsu.ldq_4_bits_debug_wb_data = 64'b0000000000000000000000000000000000000000000000000000000010100000;
    UUT.wrapper.uut.lsu.ldq_4_bits_executed = 1'b1;
    UUT.wrapper.uut.lsu.ldq_4_bits_forward_std_val = 1'b0;
    UUT.wrapper.uut.lsu.ldq_4_bits_forward_stq_idx = 4'b0001;
    UUT.wrapper.uut.lsu.ldq_4_bits_observed = 1'b0;
    UUT.wrapper.uut.lsu.ldq_4_bits_order_fail = 1'b0;
    UUT.wrapper.uut.lsu.ldq_4_bits_st_dep_mask = 16'b0000000000000000;
    UUT.wrapper.uut.lsu.ldq_4_bits_succeeded = 1'b0;
    UUT.wrapper.uut.lsu.ldq_4_bits_uop_br_mask = 12'b000000010000;
    UUT.wrapper.uut.lsu.ldq_4_bits_uop_dst_rtype = 2'b00;
    UUT.wrapper.uut.lsu.ldq_4_bits_uop_is_amo = 1'b0;
    UUT.wrapper.uut.lsu.ldq_4_bits_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_4_bits_uop_mem_cmd = 5'b00000;
    UUT.wrapper.uut.lsu.ldq_4_bits_uop_mem_signed = 1'b1;
    UUT.wrapper.uut.lsu.ldq_4_bits_uop_mem_size = 2'b10;
    UUT.wrapper.uut.lsu.ldq_4_bits_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.lsu.ldq_4_bits_uop_rob_idx = 6'b001000;
    UUT.wrapper.uut.lsu.ldq_4_bits_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_4_bits_uop_uses_ldq = 1'b1;
    UUT.wrapper.uut.lsu.ldq_4_bits_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.lsu.ldq_4_bits_youngest_stq_idx = 4'b1011;
    UUT.wrapper.uut.lsu.ldq_4_valid = 1'b1;
    UUT.wrapper.uut.lsu.ldq_5_bits_addr_bits = 40'b0001100111111111111111111111100111011111;
    UUT.wrapper.uut.lsu.ldq_5_bits_addr_is_uncacheable = 1'b1;
    UUT.wrapper.uut.lsu.ldq_5_bits_addr_is_virtual = 1'b1;
    UUT.wrapper.uut.lsu.ldq_5_bits_addr_valid = 1'b1;
    UUT.wrapper.uut.lsu.ldq_5_bits_debug_wb_data = 64'b1111111111111111111111111111111111111111111111111111111111111111;
    UUT.wrapper.uut.lsu.ldq_5_bits_executed = 1'b1;
    UUT.wrapper.uut.lsu.ldq_5_bits_forward_std_val = 1'b0;
    UUT.wrapper.uut.lsu.ldq_5_bits_forward_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_5_bits_observed = 1'b0;
    UUT.wrapper.uut.lsu.ldq_5_bits_order_fail = 1'b0;
    UUT.wrapper.uut.lsu.ldq_5_bits_st_dep_mask = 16'b0000000000000000;
    UUT.wrapper.uut.lsu.ldq_5_bits_succeeded = 1'b0;
    UUT.wrapper.uut.lsu.ldq_5_bits_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.lsu.ldq_5_bits_uop_dst_rtype = 2'b10;
    UUT.wrapper.uut.lsu.ldq_5_bits_uop_is_amo = 1'b0;
    UUT.wrapper.uut.lsu.ldq_5_bits_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_5_bits_uop_mem_cmd = 5'b00000;
    UUT.wrapper.uut.lsu.ldq_5_bits_uop_mem_signed = 1'b1;
    UUT.wrapper.uut.lsu.ldq_5_bits_uop_mem_size = 2'b11;
    UUT.wrapper.uut.lsu.ldq_5_bits_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.lsu.ldq_5_bits_uop_rob_idx = 6'b001000;
    UUT.wrapper.uut.lsu.ldq_5_bits_uop_stq_idx = 4'b0001;
    UUT.wrapper.uut.lsu.ldq_5_bits_uop_uses_ldq = 1'b1;
    UUT.wrapper.uut.lsu.ldq_5_bits_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.lsu.ldq_5_bits_youngest_stq_idx = 4'b1110;
    UUT.wrapper.uut.lsu.ldq_5_valid = 1'b1;
    UUT.wrapper.uut.lsu.ldq_6_bits_addr_bits = 40'b0001100110011001100110011001000111011111;
    UUT.wrapper.uut.lsu.ldq_6_bits_addr_is_uncacheable = 1'b1;
    UUT.wrapper.uut.lsu.ldq_6_bits_addr_is_virtual = 1'b1;
    UUT.wrapper.uut.lsu.ldq_6_bits_addr_valid = 1'b1;
    UUT.wrapper.uut.lsu.ldq_6_bits_debug_wb_data = 64'b1111111111111111111111111111111111111111111111111111111111111111;
    UUT.wrapper.uut.lsu.ldq_6_bits_executed = 1'b1;
    UUT.wrapper.uut.lsu.ldq_6_bits_forward_std_val = 1'b0;
    UUT.wrapper.uut.lsu.ldq_6_bits_forward_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_6_bits_observed = 1'b0;
    UUT.wrapper.uut.lsu.ldq_6_bits_order_fail = 1'b0;
    UUT.wrapper.uut.lsu.ldq_6_bits_st_dep_mask = 16'b0000000000000001;
    UUT.wrapper.uut.lsu.ldq_6_bits_succeeded = 1'b0;
    UUT.wrapper.uut.lsu.ldq_6_bits_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.lsu.ldq_6_bits_uop_dst_rtype = 2'b10;
    UUT.wrapper.uut.lsu.ldq_6_bits_uop_is_amo = 1'b0;
    UUT.wrapper.uut.lsu.ldq_6_bits_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_6_bits_uop_mem_cmd = 5'b00000;
    UUT.wrapper.uut.lsu.ldq_6_bits_uop_mem_signed = 1'b1;
    UUT.wrapper.uut.lsu.ldq_6_bits_uop_mem_size = 2'b11;
    UUT.wrapper.uut.lsu.ldq_6_bits_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.lsu.ldq_6_bits_uop_rob_idx = 6'b100001;
    UUT.wrapper.uut.lsu.ldq_6_bits_uop_stq_idx = 4'b0001;
    UUT.wrapper.uut.lsu.ldq_6_bits_uop_uses_ldq = 1'b1;
    UUT.wrapper.uut.lsu.ldq_6_bits_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.lsu.ldq_6_bits_youngest_stq_idx = 4'b0001;
    UUT.wrapper.uut.lsu.ldq_6_valid = 1'b1;
    UUT.wrapper.uut.lsu.ldq_7_bits_addr_bits = 40'b0001100111111111111111111111100111011111;
    UUT.wrapper.uut.lsu.ldq_7_bits_addr_is_uncacheable = 1'b1;
    UUT.wrapper.uut.lsu.ldq_7_bits_addr_is_virtual = 1'b1;
    UUT.wrapper.uut.lsu.ldq_7_bits_addr_valid = 1'b1;
    UUT.wrapper.uut.lsu.ldq_7_bits_debug_wb_data = 64'b1111111111111111111111111111111111111111111111111111111111111111;
    UUT.wrapper.uut.lsu.ldq_7_bits_executed = 1'b1;
    UUT.wrapper.uut.lsu.ldq_7_bits_forward_std_val = 1'b1;
    UUT.wrapper.uut.lsu.ldq_7_bits_forward_stq_idx = 4'b1100;
    UUT.wrapper.uut.lsu.ldq_7_bits_observed = 1'b0;
    UUT.wrapper.uut.lsu.ldq_7_bits_order_fail = 1'b1;
    UUT.wrapper.uut.lsu.ldq_7_bits_st_dep_mask = 16'b1110111111111110;
    UUT.wrapper.uut.lsu.ldq_7_bits_succeeded = 1'b1;
    UUT.wrapper.uut.lsu.ldq_7_bits_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.lsu.ldq_7_bits_uop_dst_rtype = 2'b11;
    UUT.wrapper.uut.lsu.ldq_7_bits_uop_is_amo = 1'b1;
    UUT.wrapper.uut.lsu.ldq_7_bits_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_7_bits_uop_mem_cmd = 5'b00000;
    UUT.wrapper.uut.lsu.ldq_7_bits_uop_mem_signed = 1'b1;
    UUT.wrapper.uut.lsu.ldq_7_bits_uop_mem_size = 2'b11;
    UUT.wrapper.uut.lsu.ldq_7_bits_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.lsu.ldq_7_bits_uop_rob_idx = 6'b000000;
    UUT.wrapper.uut.lsu.ldq_7_bits_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_7_bits_uop_uses_ldq = 1'b1;
    UUT.wrapper.uut.lsu.ldq_7_bits_uop_uses_stq = 1'b1;
    UUT.wrapper.uut.lsu.ldq_7_bits_youngest_stq_idx = 4'b1001;
    UUT.wrapper.uut.lsu.ldq_7_valid = 1'b1;
    UUT.wrapper.uut.lsu.ldq_8_bits_addr_bits = 40'b0001100111111111111111111111100111011111;
    UUT.wrapper.uut.lsu.ldq_8_bits_addr_is_uncacheable = 1'b1;
    UUT.wrapper.uut.lsu.ldq_8_bits_addr_is_virtual = 1'b1;
    UUT.wrapper.uut.lsu.ldq_8_bits_addr_valid = 1'b1;
    UUT.wrapper.uut.lsu.ldq_8_bits_debug_wb_data = 64'b1111111111111111111111111111111111111111111111111111111111111111;
    UUT.wrapper.uut.lsu.ldq_8_bits_executed = 1'b1;
    UUT.wrapper.uut.lsu.ldq_8_bits_forward_std_val = 1'b1;
    UUT.wrapper.uut.lsu.ldq_8_bits_forward_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_8_bits_observed = 1'b0;
    UUT.wrapper.uut.lsu.ldq_8_bits_order_fail = 1'b1;
    UUT.wrapper.uut.lsu.ldq_8_bits_st_dep_mask = 16'b1111111111111100;
    UUT.wrapper.uut.lsu.ldq_8_bits_succeeded = 1'b1;
    UUT.wrapper.uut.lsu.ldq_8_bits_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.lsu.ldq_8_bits_uop_dst_rtype = 2'b11;
    UUT.wrapper.uut.lsu.ldq_8_bits_uop_is_amo = 1'b1;
    UUT.wrapper.uut.lsu.ldq_8_bits_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_8_bits_uop_mem_cmd = 5'b00000;
    UUT.wrapper.uut.lsu.ldq_8_bits_uop_mem_signed = 1'b1;
    UUT.wrapper.uut.lsu.ldq_8_bits_uop_mem_size = 2'b11;
    UUT.wrapper.uut.lsu.ldq_8_bits_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.lsu.ldq_8_bits_uop_rob_idx = 6'b000000;
    UUT.wrapper.uut.lsu.ldq_8_bits_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_8_bits_uop_uses_ldq = 1'b1;
    UUT.wrapper.uut.lsu.ldq_8_bits_uop_uses_stq = 1'b1;
    UUT.wrapper.uut.lsu.ldq_8_bits_youngest_stq_idx = 4'b0111;
    UUT.wrapper.uut.lsu.ldq_8_valid = 1'b1;
    UUT.wrapper.uut.lsu.ldq_9_bits_addr_bits = 40'b0001100111111111111111111111100111011111;
    UUT.wrapper.uut.lsu.ldq_9_bits_addr_is_uncacheable = 1'b1;
    UUT.wrapper.uut.lsu.ldq_9_bits_addr_is_virtual = 1'b1;
    UUT.wrapper.uut.lsu.ldq_9_bits_addr_valid = 1'b1;
    UUT.wrapper.uut.lsu.ldq_9_bits_debug_wb_data = 64'b1111111111111111111111111111111111111111111111111111111111111111;
    UUT.wrapper.uut.lsu.ldq_9_bits_executed = 1'b1;
    UUT.wrapper.uut.lsu.ldq_9_bits_forward_std_val = 1'b1;
    UUT.wrapper.uut.lsu.ldq_9_bits_forward_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_9_bits_observed = 1'b0;
    UUT.wrapper.uut.lsu.ldq_9_bits_order_fail = 1'b1;
    UUT.wrapper.uut.lsu.ldq_9_bits_st_dep_mask = 16'b1111111111111110;
    UUT.wrapper.uut.lsu.ldq_9_bits_succeeded = 1'b1;
    UUT.wrapper.uut.lsu.ldq_9_bits_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.lsu.ldq_9_bits_uop_dst_rtype = 2'b11;
    UUT.wrapper.uut.lsu.ldq_9_bits_uop_is_amo = 1'b1;
    UUT.wrapper.uut.lsu.ldq_9_bits_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_9_bits_uop_mem_cmd = 5'b00000;
    UUT.wrapper.uut.lsu.ldq_9_bits_uop_mem_signed = 1'b1;
    UUT.wrapper.uut.lsu.ldq_9_bits_uop_mem_size = 2'b11;
    UUT.wrapper.uut.lsu.ldq_9_bits_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.lsu.ldq_9_bits_uop_rob_idx = 6'b000000;
    UUT.wrapper.uut.lsu.ldq_9_bits_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_9_bits_uop_uses_ldq = 1'b1;
    UUT.wrapper.uut.lsu.ldq_9_bits_uop_uses_stq = 1'b1;
    UUT.wrapper.uut.lsu.ldq_9_bits_youngest_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.ldq_9_valid = 1'b1;
    UUT.wrapper.uut.lsu.ldq_head = 4'b1111;
    UUT.wrapper.uut.lsu.ldq_retry_idx = 4'b1111;
    UUT.wrapper.uut.lsu.ldq_tail = 4'b0011;
    UUT.wrapper.uut.lsu.ldq_wakeup_idx = 4'b0010;
    UUT.wrapper.uut.lsu.live_store_mask = 16'b0000000000000001;
    UUT.wrapper.uut.lsu.mem_incoming_uop_0_br_mask = 12'b000000000000;
    UUT.wrapper.uut.lsu.mem_incoming_uop_0_fp_val = 1'b0;
    UUT.wrapper.uut.lsu.mem_incoming_uop_0_ldq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.mem_incoming_uop_0_pdst = 7'b0000000;
    UUT.wrapper.uut.lsu.mem_incoming_uop_0_rob_idx = 6'b000000;
    UUT.wrapper.uut.lsu.mem_incoming_uop_0_stq_idx = 4'b0101;
    UUT.wrapper.uut.lsu.mem_ldq_incoming_e_0_bits_st_dep_mask = 16'b1111111111111111;
    UUT.wrapper.uut.lsu.mem_ldq_incoming_e_0_bits_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.lsu.mem_ldq_incoming_e_0_bits_uop_mem_size = 2'b00;
    UUT.wrapper.uut.lsu.mem_ldq_incoming_e_0_bits_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.mem_ldq_retry_e_bits_st_dep_mask = 16'b1111111111111111;
    UUT.wrapper.uut.lsu.mem_ldq_retry_e_bits_uop_br_mask = 12'b111111111111;
    UUT.wrapper.uut.lsu.mem_ldq_retry_e_bits_uop_mem_size = 2'b11;
    UUT.wrapper.uut.lsu.mem_ldq_retry_e_bits_uop_stq_idx = 4'b1111;
    UUT.wrapper.uut.lsu.mem_ldq_wakeup_e_bits_st_dep_mask = 16'b0000000000000000;
    UUT.wrapper.uut.lsu.mem_ldq_wakeup_e_bits_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.lsu.mem_ldq_wakeup_e_bits_uop_mem_size = 2'b00;
    UUT.wrapper.uut.lsu.mem_ldq_wakeup_e_bits_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.mem_paddr_0 = 40'b1111111100000000000000000000000000000010;
    UUT.wrapper.uut.lsu.mem_stq_incoming_e_0_bits_addr_is_virtual = 1'b0;
    UUT.wrapper.uut.lsu.mem_stq_incoming_e_0_bits_addr_valid = 1'b0;
    UUT.wrapper.uut.lsu.mem_stq_incoming_e_0_bits_data_valid = 1'b0;
    UUT.wrapper.uut.lsu.mem_stq_incoming_e_0_bits_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.lsu.mem_stq_incoming_e_0_bits_uop_is_amo = 1'b0;
    UUT.wrapper.uut.lsu.mem_stq_incoming_e_0_bits_uop_mem_size = 2'b00;
    UUT.wrapper.uut.lsu.mem_stq_incoming_e_0_bits_uop_rob_idx = 6'b000000;
    UUT.wrapper.uut.lsu.mem_stq_incoming_e_0_bits_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.mem_stq_incoming_e_0_valid = 1'b0;
    UUT.wrapper.uut.lsu.mem_stq_retry_e_bits_data_valid = 1'b0;
    UUT.wrapper.uut.lsu.mem_stq_retry_e_bits_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.lsu.mem_stq_retry_e_bits_uop_is_amo = 1'b0;
    UUT.wrapper.uut.lsu.mem_stq_retry_e_bits_uop_mem_size = 2'b01;
    UUT.wrapper.uut.lsu.mem_stq_retry_e_bits_uop_rob_idx = 6'b000000;
    UUT.wrapper.uut.lsu.mem_stq_retry_e_bits_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.mem_stq_retry_e_valid = 1'b0;
    UUT.wrapper.uut.lsu.mem_tlb_miss_0 = 1'b1;
    UUT.wrapper.uut.lsu.mem_tlb_uncacheable_0 = 1'b0;
    UUT.wrapper.uut.lsu.mem_xcpt_causes_0 = 4'b0000;
    UUT.wrapper.uut.lsu.mem_xcpt_uops_0_br_mask = 12'b000000000000;
    UUT.wrapper.uut.lsu.mem_xcpt_uops_0_rob_idx = 6'b000000;
    UUT.wrapper.uut.lsu.mem_xcpt_uops_0_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.mem_xcpt_uops_0_uses_ldq = 1'b0;
    UUT.wrapper.uut.lsu.mem_xcpt_vaddrs_0 = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.lsu.mem_xcpt_valids_0 = 1'b1;
    UUT.wrapper.uut.lsu.older_nacked_REG = 1'b0;
    UUT.wrapper.uut.lsu.older_nacked_REG_1 = 1'b1;
    UUT.wrapper.uut.lsu.older_nacked_REG_10 = 1'b1;
    UUT.wrapper.uut.lsu.older_nacked_REG_11 = 1'b0;
    UUT.wrapper.uut.lsu.older_nacked_REG_12 = 1'b1;
    UUT.wrapper.uut.lsu.older_nacked_REG_13 = 1'b1;
    UUT.wrapper.uut.lsu.older_nacked_REG_14 = 1'b1;
    UUT.wrapper.uut.lsu.older_nacked_REG_15 = 1'b1;
    UUT.wrapper.uut.lsu.older_nacked_REG_2 = 1'b1;
    UUT.wrapper.uut.lsu.older_nacked_REG_3 = 1'b1;
    UUT.wrapper.uut.lsu.older_nacked_REG_4 = 1'b1;
    UUT.wrapper.uut.lsu.older_nacked_REG_5 = 1'b1;
    UUT.wrapper.uut.lsu.older_nacked_REG_6 = 1'b1;
    UUT.wrapper.uut.lsu.older_nacked_REG_7 = 1'b1;
    UUT.wrapper.uut.lsu.older_nacked_REG_8 = 1'b1;
    UUT.wrapper.uut.lsu.older_nacked_REG_9 = 1'b1;
    UUT.wrapper.uut.lsu.p1_block_load_mask_0 = 1'b1;
    UUT.wrapper.uut.lsu.p1_block_load_mask_1 = 1'b1;
    UUT.wrapper.uut.lsu.p1_block_load_mask_10 = 1'b1;
    UUT.wrapper.uut.lsu.p1_block_load_mask_11 = 1'b1;
    UUT.wrapper.uut.lsu.p1_block_load_mask_12 = 1'b1;
    UUT.wrapper.uut.lsu.p1_block_load_mask_13 = 1'b1;
    UUT.wrapper.uut.lsu.p1_block_load_mask_14 = 1'b1;
    UUT.wrapper.uut.lsu.p1_block_load_mask_15 = 1'b0;
    UUT.wrapper.uut.lsu.p1_block_load_mask_2 = 1'b1;
    UUT.wrapper.uut.lsu.p1_block_load_mask_3 = 1'b1;
    UUT.wrapper.uut.lsu.p1_block_load_mask_4 = 1'b1;
    UUT.wrapper.uut.lsu.p1_block_load_mask_5 = 1'b0;
    UUT.wrapper.uut.lsu.p1_block_load_mask_6 = 1'b1;
    UUT.wrapper.uut.lsu.p1_block_load_mask_7 = 1'b1;
    UUT.wrapper.uut.lsu.p1_block_load_mask_8 = 1'b1;
    UUT.wrapper.uut.lsu.p1_block_load_mask_9 = 1'b1;
    UUT.wrapper.uut.lsu.p2_block_load_mask_0 = 1'b1;
    UUT.wrapper.uut.lsu.p2_block_load_mask_1 = 1'b1;
    UUT.wrapper.uut.lsu.p2_block_load_mask_10 = 1'b1;
    UUT.wrapper.uut.lsu.p2_block_load_mask_11 = 1'b1;
    UUT.wrapper.uut.lsu.p2_block_load_mask_12 = 1'b1;
    UUT.wrapper.uut.lsu.p2_block_load_mask_13 = 1'b1;
    UUT.wrapper.uut.lsu.p2_block_load_mask_14 = 1'b1;
    UUT.wrapper.uut.lsu.p2_block_load_mask_15 = 1'b0;
    UUT.wrapper.uut.lsu.p2_block_load_mask_2 = 1'b1;
    UUT.wrapper.uut.lsu.p2_block_load_mask_3 = 1'b1;
    UUT.wrapper.uut.lsu.p2_block_load_mask_4 = 1'b1;
    UUT.wrapper.uut.lsu.p2_block_load_mask_5 = 1'b0;
    UUT.wrapper.uut.lsu.p2_block_load_mask_6 = 1'b1;
    UUT.wrapper.uut.lsu.p2_block_load_mask_7 = 1'b1;
    UUT.wrapper.uut.lsu.p2_block_load_mask_8 = 1'b1;
    UUT.wrapper.uut.lsu.p2_block_load_mask_9 = 1'b1;
    UUT.wrapper.uut.lsu.r_xcpt_badvaddr = 40'b0000000000000000000000000000000000000000;
    UUT.wrapper.uut.lsu.r_xcpt_cause = 5'b00000;
    UUT.wrapper.uut.lsu.r_xcpt_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.lsu.r_xcpt_uop_rob_idx = 6'b000000;
    UUT.wrapper.uut.lsu.r_xcpt_valid = 1'b0;
    UUT.wrapper.uut.lsu.s1_executing_loads_0 = 1'b1;
    UUT.wrapper.uut.lsu.s1_executing_loads_1 = 1'b1;
    UUT.wrapper.uut.lsu.s1_executing_loads_10 = 1'b0;
    UUT.wrapper.uut.lsu.s1_executing_loads_11 = 1'b0;
    UUT.wrapper.uut.lsu.s1_executing_loads_12 = 1'b0;
    UUT.wrapper.uut.lsu.s1_executing_loads_13 = 1'b0;
    UUT.wrapper.uut.lsu.s1_executing_loads_14 = 1'b0;
    UUT.wrapper.uut.lsu.s1_executing_loads_15 = 1'b0;
    UUT.wrapper.uut.lsu.s1_executing_loads_2 = 1'b0;
    UUT.wrapper.uut.lsu.s1_executing_loads_3 = 1'b0;
    UUT.wrapper.uut.lsu.s1_executing_loads_4 = 1'b0;
    UUT.wrapper.uut.lsu.s1_executing_loads_5 = 1'b1;
    UUT.wrapper.uut.lsu.s1_executing_loads_6 = 1'b0;
    UUT.wrapper.uut.lsu.s1_executing_loads_7 = 1'b1;
    UUT.wrapper.uut.lsu.s1_executing_loads_8 = 1'b0;
    UUT.wrapper.uut.lsu.s1_executing_loads_9 = 1'b0;
    UUT.wrapper.uut.lsu.spec_ld_succeed_REG = 1'b1;
    UUT.wrapper.uut.lsu.spec_ld_succeed_REG_1 = 4'b1000;
    UUT.wrapper.uut.lsu.store_blocked_counter = 4'b1110;
    UUT.wrapper.uut.lsu.stq_0_bits_addr_bits = 40'b0000000001000110000000000111100000000000;
    UUT.wrapper.uut.lsu.stq_0_bits_addr_is_virtual = 1'b0;
    UUT.wrapper.uut.lsu.stq_0_bits_addr_valid = 1'b1;
    UUT.wrapper.uut.lsu.stq_0_bits_committed = 1'b1;
    UUT.wrapper.uut.lsu.stq_0_bits_data_bits = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.lsu.stq_0_bits_data_valid = 1'b0;
    UUT.wrapper.uut.lsu.stq_0_bits_debug_wb_data = 64'b0000000000000000000000000000000000000000000000000000000000001000;
    UUT.wrapper.uut.lsu.stq_0_bits_succeeded = 1'b1;
    UUT.wrapper.uut.lsu.stq_0_bits_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.lsu.stq_0_bits_uop_dst_rtype = 2'b00;
    UUT.wrapper.uut.lsu.stq_0_bits_uop_exception = 1'b0;
    UUT.wrapper.uut.lsu.stq_0_bits_uop_is_amo = 1'b1;
    UUT.wrapper.uut.lsu.stq_0_bits_uop_is_fence = 1'b0;
    UUT.wrapper.uut.lsu.stq_0_bits_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.stq_0_bits_uop_mem_cmd = 5'b10001;
    UUT.wrapper.uut.lsu.stq_0_bits_uop_mem_signed = 1'b0;
    UUT.wrapper.uut.lsu.stq_0_bits_uop_mem_size = 2'b00;
    UUT.wrapper.uut.lsu.stq_0_bits_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.lsu.stq_0_bits_uop_rob_idx = 6'b000001;
    UUT.wrapper.uut.lsu.stq_0_bits_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.stq_0_bits_uop_uses_ldq = 1'b0;
    UUT.wrapper.uut.lsu.stq_0_bits_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.lsu.stq_0_valid = 1'b0;
    UUT.wrapper.uut.lsu.stq_10_bits_addr_bits = 40'b0000000011111111111111111111100110011111;
    UUT.wrapper.uut.lsu.stq_10_bits_addr_is_virtual = 1'b1;
    UUT.wrapper.uut.lsu.stq_10_bits_addr_valid = 1'b1;
    UUT.wrapper.uut.lsu.stq_10_bits_committed = 1'b1;
    UUT.wrapper.uut.lsu.stq_10_bits_data_bits = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.lsu.stq_10_bits_data_valid = 1'b0;
    UUT.wrapper.uut.lsu.stq_10_bits_debug_wb_data = 64'b1111111111111111111111111111111111111111111111111111111111111111;
    UUT.wrapper.uut.lsu.stq_10_bits_succeeded = 1'b1;
    UUT.wrapper.uut.lsu.stq_10_bits_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.lsu.stq_10_bits_uop_dst_rtype = 2'b11;
    UUT.wrapper.uut.lsu.stq_10_bits_uop_exception = 1'b0;
    UUT.wrapper.uut.lsu.stq_10_bits_uop_is_amo = 1'b1;
    UUT.wrapper.uut.lsu.stq_10_bits_uop_is_fence = 1'b1;
    UUT.wrapper.uut.lsu.stq_10_bits_uop_ldq_idx = 4'b1111;
    UUT.wrapper.uut.lsu.stq_10_bits_uop_mem_cmd = 5'b11111;
    UUT.wrapper.uut.lsu.stq_10_bits_uop_mem_signed = 1'b0;
    UUT.wrapper.uut.lsu.stq_10_bits_uop_mem_size = 2'b00;
    UUT.wrapper.uut.lsu.stq_10_bits_uop_pdst = 7'b1111111;
    UUT.wrapper.uut.lsu.stq_10_bits_uop_rob_idx = 6'b111111;
    UUT.wrapper.uut.lsu.stq_10_bits_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.stq_10_bits_uop_uses_ldq = 1'b0;
    UUT.wrapper.uut.lsu.stq_10_bits_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.lsu.stq_10_valid = 1'b1;
    UUT.wrapper.uut.lsu.stq_11_bits_addr_bits = 40'b0000000011111111111111111111100110011011;
    UUT.wrapper.uut.lsu.stq_11_bits_addr_is_virtual = 1'b1;
    UUT.wrapper.uut.lsu.stq_11_bits_addr_valid = 1'b0;
    UUT.wrapper.uut.lsu.stq_11_bits_committed = 1'b1;
    UUT.wrapper.uut.lsu.stq_11_bits_data_bits = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.lsu.stq_11_bits_data_valid = 1'b1;
    UUT.wrapper.uut.lsu.stq_11_bits_debug_wb_data = 64'b1111111111111111111111111111111111111111111111111111111111111111;
    UUT.wrapper.uut.lsu.stq_11_bits_succeeded = 1'b1;
    UUT.wrapper.uut.lsu.stq_11_bits_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.lsu.stq_11_bits_uop_dst_rtype = 2'b11;
    UUT.wrapper.uut.lsu.stq_11_bits_uop_exception = 1'b1;
    UUT.wrapper.uut.lsu.stq_11_bits_uop_is_amo = 1'b1;
    UUT.wrapper.uut.lsu.stq_11_bits_uop_is_fence = 1'b1;
    UUT.wrapper.uut.lsu.stq_11_bits_uop_ldq_idx = 4'b1111;
    UUT.wrapper.uut.lsu.stq_11_bits_uop_mem_cmd = 5'b11111;
    UUT.wrapper.uut.lsu.stq_11_bits_uop_mem_signed = 1'b0;
    UUT.wrapper.uut.lsu.stq_11_bits_uop_mem_size = 2'b00;
    UUT.wrapper.uut.lsu.stq_11_bits_uop_pdst = 7'b1111111;
    UUT.wrapper.uut.lsu.stq_11_bits_uop_rob_idx = 6'b111111;
    UUT.wrapper.uut.lsu.stq_11_bits_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.stq_11_bits_uop_uses_ldq = 1'b0;
    UUT.wrapper.uut.lsu.stq_11_bits_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.lsu.stq_11_valid = 1'b1;
    UUT.wrapper.uut.lsu.stq_12_bits_addr_bits = 40'b1110011011111111111111111111000000011111;
    UUT.wrapper.uut.lsu.stq_12_bits_addr_is_virtual = 1'b1;
    UUT.wrapper.uut.lsu.stq_12_bits_addr_valid = 1'b0;
    UUT.wrapper.uut.lsu.stq_12_bits_committed = 1'b1;
    UUT.wrapper.uut.lsu.stq_12_bits_data_bits = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.lsu.stq_12_bits_data_valid = 1'b0;
    UUT.wrapper.uut.lsu.stq_12_bits_debug_wb_data = 64'b1111111111111111111111111111111111111111111111111111111111111111;
    UUT.wrapper.uut.lsu.stq_12_bits_succeeded = 1'b1;
    UUT.wrapper.uut.lsu.stq_12_bits_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.lsu.stq_12_bits_uop_dst_rtype = 2'b11;
    UUT.wrapper.uut.lsu.stq_12_bits_uop_exception = 1'b1;
    UUT.wrapper.uut.lsu.stq_12_bits_uop_is_amo = 1'b0;
    UUT.wrapper.uut.lsu.stq_12_bits_uop_is_fence = 1'b1;
    UUT.wrapper.uut.lsu.stq_12_bits_uop_ldq_idx = 4'b1111;
    UUT.wrapper.uut.lsu.stq_12_bits_uop_mem_cmd = 5'b11111;
    UUT.wrapper.uut.lsu.stq_12_bits_uop_mem_signed = 1'b0;
    UUT.wrapper.uut.lsu.stq_12_bits_uop_mem_size = 2'b00;
    UUT.wrapper.uut.lsu.stq_12_bits_uop_pdst = 7'b1111111;
    UUT.wrapper.uut.lsu.stq_12_bits_uop_rob_idx = 6'b111111;
    UUT.wrapper.uut.lsu.stq_12_bits_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.stq_12_bits_uop_uses_ldq = 1'b0;
    UUT.wrapper.uut.lsu.stq_12_bits_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.lsu.stq_12_valid = 1'b1;
    UUT.wrapper.uut.lsu.stq_13_bits_addr_bits = 40'b0000000011111111111111111111100110011111;
    UUT.wrapper.uut.lsu.stq_13_bits_addr_is_virtual = 1'b1;
    UUT.wrapper.uut.lsu.stq_13_bits_addr_valid = 1'b0;
    UUT.wrapper.uut.lsu.stq_13_bits_committed = 1'b1;
    UUT.wrapper.uut.lsu.stq_13_bits_data_bits = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.lsu.stq_13_bits_data_valid = 1'b1;
    UUT.wrapper.uut.lsu.stq_13_bits_debug_wb_data = 64'b1111111111111111111111111111111111111111111111111111111111111111;
    UUT.wrapper.uut.lsu.stq_13_bits_succeeded = 1'b1;
    UUT.wrapper.uut.lsu.stq_13_bits_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.lsu.stq_13_bits_uop_dst_rtype = 2'b11;
    UUT.wrapper.uut.lsu.stq_13_bits_uop_exception = 1'b1;
    UUT.wrapper.uut.lsu.stq_13_bits_uop_is_amo = 1'b0;
    UUT.wrapper.uut.lsu.stq_13_bits_uop_is_fence = 1'b1;
    UUT.wrapper.uut.lsu.stq_13_bits_uop_ldq_idx = 4'b1111;
    UUT.wrapper.uut.lsu.stq_13_bits_uop_mem_cmd = 5'b11111;
    UUT.wrapper.uut.lsu.stq_13_bits_uop_mem_signed = 1'b0;
    UUT.wrapper.uut.lsu.stq_13_bits_uop_mem_size = 2'b00;
    UUT.wrapper.uut.lsu.stq_13_bits_uop_pdst = 7'b1111111;
    UUT.wrapper.uut.lsu.stq_13_bits_uop_rob_idx = 6'b111111;
    UUT.wrapper.uut.lsu.stq_13_bits_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.stq_13_bits_uop_uses_ldq = 1'b0;
    UUT.wrapper.uut.lsu.stq_13_bits_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.lsu.stq_13_valid = 1'b1;
    UUT.wrapper.uut.lsu.stq_14_bits_addr_bits = 40'b1110010011111111111111111111100110011111;
    UUT.wrapper.uut.lsu.stq_14_bits_addr_is_virtual = 1'b1;
    UUT.wrapper.uut.lsu.stq_14_bits_addr_valid = 1'b0;
    UUT.wrapper.uut.lsu.stq_14_bits_committed = 1'b1;
    UUT.wrapper.uut.lsu.stq_14_bits_data_bits = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.lsu.stq_14_bits_data_valid = 1'b0;
    UUT.wrapper.uut.lsu.stq_14_bits_debug_wb_data = 64'b1111111111111111111111111111111111111111111111111111111111111111;
    UUT.wrapper.uut.lsu.stq_14_bits_succeeded = 1'b1;
    UUT.wrapper.uut.lsu.stq_14_bits_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.lsu.stq_14_bits_uop_dst_rtype = 2'b11;
    UUT.wrapper.uut.lsu.stq_14_bits_uop_exception = 1'b1;
    UUT.wrapper.uut.lsu.stq_14_bits_uop_is_amo = 1'b1;
    UUT.wrapper.uut.lsu.stq_14_bits_uop_is_fence = 1'b1;
    UUT.wrapper.uut.lsu.stq_14_bits_uop_ldq_idx = 4'b1111;
    UUT.wrapper.uut.lsu.stq_14_bits_uop_mem_cmd = 5'b10001;
    UUT.wrapper.uut.lsu.stq_14_bits_uop_mem_signed = 1'b0;
    UUT.wrapper.uut.lsu.stq_14_bits_uop_mem_size = 2'b00;
    UUT.wrapper.uut.lsu.stq_14_bits_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.lsu.stq_14_bits_uop_rob_idx = 6'b111111;
    UUT.wrapper.uut.lsu.stq_14_bits_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.stq_14_bits_uop_uses_ldq = 1'b0;
    UUT.wrapper.uut.lsu.stq_14_bits_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.lsu.stq_14_valid = 1'b1;
    UUT.wrapper.uut.lsu.stq_15_bits_addr_bits = 40'b1111111111110111111111111111100110011111;
    UUT.wrapper.uut.lsu.stq_15_bits_addr_is_virtual = 1'b1;
    UUT.wrapper.uut.lsu.stq_15_bits_addr_valid = 1'b1;
    UUT.wrapper.uut.lsu.stq_15_bits_committed = 1'b1;
    UUT.wrapper.uut.lsu.stq_15_bits_data_bits = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.lsu.stq_15_bits_data_valid = 1'b1;
    UUT.wrapper.uut.lsu.stq_15_bits_debug_wb_data = 64'b1111111111111111111111111111111110000000000000001000000010000000;
    UUT.wrapper.uut.lsu.stq_15_bits_succeeded = 1'b1;
    UUT.wrapper.uut.lsu.stq_15_bits_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.lsu.stq_15_bits_uop_dst_rtype = 2'b11;
    UUT.wrapper.uut.lsu.stq_15_bits_uop_exception = 1'b0;
    UUT.wrapper.uut.lsu.stq_15_bits_uop_is_amo = 1'b1;
    UUT.wrapper.uut.lsu.stq_15_bits_uop_is_fence = 1'b1;
    UUT.wrapper.uut.lsu.stq_15_bits_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.stq_15_bits_uop_mem_cmd = 5'b10001;
    UUT.wrapper.uut.lsu.stq_15_bits_uop_mem_signed = 1'b0;
    UUT.wrapper.uut.lsu.stq_15_bits_uop_mem_size = 2'b00;
    UUT.wrapper.uut.lsu.stq_15_bits_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.lsu.stq_15_bits_uop_rob_idx = 6'b000101;
    UUT.wrapper.uut.lsu.stq_15_bits_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.stq_15_bits_uop_uses_ldq = 1'b0;
    UUT.wrapper.uut.lsu.stq_15_bits_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.lsu.stq_15_valid = 1'b1;
    UUT.wrapper.uut.lsu.stq_1_bits_addr_bits = 40'b0000000000010000000000000000000000010000;
    UUT.wrapper.uut.lsu.stq_1_bits_addr_is_virtual = 1'b0;
    UUT.wrapper.uut.lsu.stq_1_bits_addr_valid = 1'b1;
    UUT.wrapper.uut.lsu.stq_1_bits_committed = 1'b0;
    UUT.wrapper.uut.lsu.stq_1_bits_data_bits = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.lsu.stq_1_bits_data_valid = 1'b0;
    UUT.wrapper.uut.lsu.stq_1_bits_debug_wb_data = 64'b1111111111111111111111111111111111111111111111111111111111111110;
    UUT.wrapper.uut.lsu.stq_1_bits_succeeded = 1'b0;
    UUT.wrapper.uut.lsu.stq_1_bits_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.lsu.stq_1_bits_uop_dst_rtype = 2'b00;
    UUT.wrapper.uut.lsu.stq_1_bits_uop_exception = 1'b0;
    UUT.wrapper.uut.lsu.stq_1_bits_uop_is_amo = 1'b1;
    UUT.wrapper.uut.lsu.stq_1_bits_uop_is_fence = 1'b1;
    UUT.wrapper.uut.lsu.stq_1_bits_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.stq_1_bits_uop_mem_cmd = 5'b00000;
    UUT.wrapper.uut.lsu.stq_1_bits_uop_mem_signed = 1'b0;
    UUT.wrapper.uut.lsu.stq_1_bits_uop_mem_size = 2'b00;
    UUT.wrapper.uut.lsu.stq_1_bits_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.lsu.stq_1_bits_uop_rob_idx = 6'b000000;
    UUT.wrapper.uut.lsu.stq_1_bits_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.stq_1_bits_uop_uses_ldq = 1'b0;
    UUT.wrapper.uut.lsu.stq_1_bits_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.lsu.stq_1_valid = 1'b1;
    UUT.wrapper.uut.lsu.stq_2_bits_addr_bits = 40'b0000000011100111111111111111100100001011;
    UUT.wrapper.uut.lsu.stq_2_bits_addr_is_virtual = 1'b1;
    UUT.wrapper.uut.lsu.stq_2_bits_addr_valid = 1'b0;
    UUT.wrapper.uut.lsu.stq_2_bits_committed = 1'b0;
    UUT.wrapper.uut.lsu.stq_2_bits_data_bits = 64'b0000000000000000000000011000000110000000000000001000000000100000;
    UUT.wrapper.uut.lsu.stq_2_bits_data_valid = 1'b1;
    UUT.wrapper.uut.lsu.stq_2_bits_debug_wb_data = 64'b1111111111111111111111111111111111111111111111111111111111111111;
    UUT.wrapper.uut.lsu.stq_2_bits_succeeded = 1'b0;
    UUT.wrapper.uut.lsu.stq_2_bits_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.lsu.stq_2_bits_uop_dst_rtype = 2'b11;
    UUT.wrapper.uut.lsu.stq_2_bits_uop_exception = 1'b1;
    UUT.wrapper.uut.lsu.stq_2_bits_uop_is_amo = 1'b1;
    UUT.wrapper.uut.lsu.stq_2_bits_uop_is_fence = 1'b1;
    UUT.wrapper.uut.lsu.stq_2_bits_uop_ldq_idx = 4'b1111;
    UUT.wrapper.uut.lsu.stq_2_bits_uop_mem_cmd = 5'b11111;
    UUT.wrapper.uut.lsu.stq_2_bits_uop_mem_signed = 1'b0;
    UUT.wrapper.uut.lsu.stq_2_bits_uop_mem_size = 2'b10;
    UUT.wrapper.uut.lsu.stq_2_bits_uop_pdst = 7'b1111111;
    UUT.wrapper.uut.lsu.stq_2_bits_uop_rob_idx = 6'b111111;
    UUT.wrapper.uut.lsu.stq_2_bits_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.stq_2_bits_uop_uses_ldq = 1'b0;
    UUT.wrapper.uut.lsu.stq_2_bits_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.lsu.stq_2_valid = 1'b1;
    UUT.wrapper.uut.lsu.stq_3_bits_addr_bits = 40'b0000000011111111111101111111100110001111;
    UUT.wrapper.uut.lsu.stq_3_bits_addr_is_virtual = 1'b1;
    UUT.wrapper.uut.lsu.stq_3_bits_addr_valid = 1'b1;
    UUT.wrapper.uut.lsu.stq_3_bits_committed = 1'b1;
    UUT.wrapper.uut.lsu.stq_3_bits_data_bits = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.lsu.stq_3_bits_data_valid = 1'b1;
    UUT.wrapper.uut.lsu.stq_3_bits_debug_wb_data = 64'b1111111111111111111111111111111111111111111111111111111111111111;
    UUT.wrapper.uut.lsu.stq_3_bits_succeeded = 1'b1;
    UUT.wrapper.uut.lsu.stq_3_bits_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.lsu.stq_3_bits_uop_dst_rtype = 2'b11;
    UUT.wrapper.uut.lsu.stq_3_bits_uop_exception = 1'b1;
    UUT.wrapper.uut.lsu.stq_3_bits_uop_is_amo = 1'b0;
    UUT.wrapper.uut.lsu.stq_3_bits_uop_is_fence = 1'b1;
    UUT.wrapper.uut.lsu.stq_3_bits_uop_ldq_idx = 4'b1111;
    UUT.wrapper.uut.lsu.stq_3_bits_uop_mem_cmd = 5'b11111;
    UUT.wrapper.uut.lsu.stq_3_bits_uop_mem_signed = 1'b0;
    UUT.wrapper.uut.lsu.stq_3_bits_uop_mem_size = 2'b10;
    UUT.wrapper.uut.lsu.stq_3_bits_uop_pdst = 7'b1111111;
    UUT.wrapper.uut.lsu.stq_3_bits_uop_rob_idx = 6'b111111;
    UUT.wrapper.uut.lsu.stq_3_bits_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.stq_3_bits_uop_uses_ldq = 1'b0;
    UUT.wrapper.uut.lsu.stq_3_bits_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.lsu.stq_3_valid = 1'b1;
    UUT.wrapper.uut.lsu.stq_4_bits_addr_bits = 40'b0000000011101111111111100110100110011011;
    UUT.wrapper.uut.lsu.stq_4_bits_addr_is_virtual = 1'b1;
    UUT.wrapper.uut.lsu.stq_4_bits_addr_valid = 1'b1;
    UUT.wrapper.uut.lsu.stq_4_bits_committed = 1'b1;
    UUT.wrapper.uut.lsu.stq_4_bits_data_bits = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.lsu.stq_4_bits_data_valid = 1'b1;
    UUT.wrapper.uut.lsu.stq_4_bits_debug_wb_data = 64'b1111111111111111111111111111111111111111111111111111111111111111;
    UUT.wrapper.uut.lsu.stq_4_bits_succeeded = 1'b1;
    UUT.wrapper.uut.lsu.stq_4_bits_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.lsu.stq_4_bits_uop_dst_rtype = 2'b11;
    UUT.wrapper.uut.lsu.stq_4_bits_uop_exception = 1'b1;
    UUT.wrapper.uut.lsu.stq_4_bits_uop_is_amo = 1'b1;
    UUT.wrapper.uut.lsu.stq_4_bits_uop_is_fence = 1'b1;
    UUT.wrapper.uut.lsu.stq_4_bits_uop_ldq_idx = 4'b1111;
    UUT.wrapper.uut.lsu.stq_4_bits_uop_mem_cmd = 5'b11111;
    UUT.wrapper.uut.lsu.stq_4_bits_uop_mem_signed = 1'b0;
    UUT.wrapper.uut.lsu.stq_4_bits_uop_mem_size = 2'b10;
    UUT.wrapper.uut.lsu.stq_4_bits_uop_pdst = 7'b1111111;
    UUT.wrapper.uut.lsu.stq_4_bits_uop_rob_idx = 6'b111111;
    UUT.wrapper.uut.lsu.stq_4_bits_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.stq_4_bits_uop_uses_ldq = 1'b0;
    UUT.wrapper.uut.lsu.stq_4_bits_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.lsu.stq_4_valid = 1'b1;
    UUT.wrapper.uut.lsu.stq_5_bits_addr_bits = 40'b0000000011111111111111111111100110011110;
    UUT.wrapper.uut.lsu.stq_5_bits_addr_is_virtual = 1'b1;
    UUT.wrapper.uut.lsu.stq_5_bits_addr_valid = 1'b0;
    UUT.wrapper.uut.lsu.stq_5_bits_committed = 1'b1;
    UUT.wrapper.uut.lsu.stq_5_bits_data_bits = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.lsu.stq_5_bits_data_valid = 1'b1;
    UUT.wrapper.uut.lsu.stq_5_bits_debug_wb_data = 64'b1111111111111111111111111111111111111111111111111111111111111111;
    UUT.wrapper.uut.lsu.stq_5_bits_succeeded = 1'b1;
    UUT.wrapper.uut.lsu.stq_5_bits_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.lsu.stq_5_bits_uop_dst_rtype = 2'b11;
    UUT.wrapper.uut.lsu.stq_5_bits_uop_exception = 1'b0;
    UUT.wrapper.uut.lsu.stq_5_bits_uop_is_amo = 1'b1;
    UUT.wrapper.uut.lsu.stq_5_bits_uop_is_fence = 1'b1;
    UUT.wrapper.uut.lsu.stq_5_bits_uop_ldq_idx = 4'b1111;
    UUT.wrapper.uut.lsu.stq_5_bits_uop_mem_cmd = 5'b11111;
    UUT.wrapper.uut.lsu.stq_5_bits_uop_mem_signed = 1'b0;
    UUT.wrapper.uut.lsu.stq_5_bits_uop_mem_size = 2'b10;
    UUT.wrapper.uut.lsu.stq_5_bits_uop_pdst = 7'b1111111;
    UUT.wrapper.uut.lsu.stq_5_bits_uop_rob_idx = 6'b111111;
    UUT.wrapper.uut.lsu.stq_5_bits_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.stq_5_bits_uop_uses_ldq = 1'b0;
    UUT.wrapper.uut.lsu.stq_5_bits_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.lsu.stq_5_valid = 1'b1;
    UUT.wrapper.uut.lsu.stq_6_bits_addr_bits = 40'b0000000011111111111111111111100100010111;
    UUT.wrapper.uut.lsu.stq_6_bits_addr_is_virtual = 1'b1;
    UUT.wrapper.uut.lsu.stq_6_bits_addr_valid = 1'b0;
    UUT.wrapper.uut.lsu.stq_6_bits_committed = 1'b1;
    UUT.wrapper.uut.lsu.stq_6_bits_data_bits = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.lsu.stq_6_bits_data_valid = 1'b0;
    UUT.wrapper.uut.lsu.stq_6_bits_debug_wb_data = 64'b1111111111111111111111111111111111111111111111111111111111111111;
    UUT.wrapper.uut.lsu.stq_6_bits_succeeded = 1'b1;
    UUT.wrapper.uut.lsu.stq_6_bits_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.lsu.stq_6_bits_uop_dst_rtype = 2'b11;
    UUT.wrapper.uut.lsu.stq_6_bits_uop_exception = 1'b1;
    UUT.wrapper.uut.lsu.stq_6_bits_uop_is_amo = 1'b1;
    UUT.wrapper.uut.lsu.stq_6_bits_uop_is_fence = 1'b1;
    UUT.wrapper.uut.lsu.stq_6_bits_uop_ldq_idx = 4'b1111;
    UUT.wrapper.uut.lsu.stq_6_bits_uop_mem_cmd = 5'b11111;
    UUT.wrapper.uut.lsu.stq_6_bits_uop_mem_signed = 1'b0;
    UUT.wrapper.uut.lsu.stq_6_bits_uop_mem_size = 2'b00;
    UUT.wrapper.uut.lsu.stq_6_bits_uop_pdst = 7'b1111111;
    UUT.wrapper.uut.lsu.stq_6_bits_uop_rob_idx = 6'b111111;
    UUT.wrapper.uut.lsu.stq_6_bits_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.stq_6_bits_uop_uses_ldq = 1'b0;
    UUT.wrapper.uut.lsu.stq_6_bits_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.lsu.stq_6_valid = 1'b1;
    UUT.wrapper.uut.lsu.stq_7_bits_addr_bits = 40'b0000000011111110111111111111100110011111;
    UUT.wrapper.uut.lsu.stq_7_bits_addr_is_virtual = 1'b1;
    UUT.wrapper.uut.lsu.stq_7_bits_addr_valid = 1'b0;
    UUT.wrapper.uut.lsu.stq_7_bits_committed = 1'b1;
    UUT.wrapper.uut.lsu.stq_7_bits_data_bits = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.lsu.stq_7_bits_data_valid = 1'b1;
    UUT.wrapper.uut.lsu.stq_7_bits_debug_wb_data = 64'b1111111111111111111111111111111111111111111111111111111111111111;
    UUT.wrapper.uut.lsu.stq_7_bits_succeeded = 1'b1;
    UUT.wrapper.uut.lsu.stq_7_bits_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.lsu.stq_7_bits_uop_dst_rtype = 2'b11;
    UUT.wrapper.uut.lsu.stq_7_bits_uop_exception = 1'b1;
    UUT.wrapper.uut.lsu.stq_7_bits_uop_is_amo = 1'b1;
    UUT.wrapper.uut.lsu.stq_7_bits_uop_is_fence = 1'b1;
    UUT.wrapper.uut.lsu.stq_7_bits_uop_ldq_idx = 4'b1111;
    UUT.wrapper.uut.lsu.stq_7_bits_uop_mem_cmd = 5'b00000;
    UUT.wrapper.uut.lsu.stq_7_bits_uop_mem_signed = 1'b0;
    UUT.wrapper.uut.lsu.stq_7_bits_uop_mem_size = 2'b00;
    UUT.wrapper.uut.lsu.stq_7_bits_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.lsu.stq_7_bits_uop_rob_idx = 6'b111111;
    UUT.wrapper.uut.lsu.stq_7_bits_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.stq_7_bits_uop_uses_ldq = 1'b0;
    UUT.wrapper.uut.lsu.stq_7_bits_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.lsu.stq_7_valid = 1'b1;
    UUT.wrapper.uut.lsu.stq_8_bits_addr_bits = 40'b0000000011111111111111111111100100011111;
    UUT.wrapper.uut.lsu.stq_8_bits_addr_is_virtual = 1'b1;
    UUT.wrapper.uut.lsu.stq_8_bits_addr_valid = 1'b0;
    UUT.wrapper.uut.lsu.stq_8_bits_committed = 1'b1;
    UUT.wrapper.uut.lsu.stq_8_bits_data_bits = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.lsu.stq_8_bits_data_valid = 1'b1;
    UUT.wrapper.uut.lsu.stq_8_bits_debug_wb_data = 64'b0000000000000000000000000000000000000000000000000000000000001000;
    UUT.wrapper.uut.lsu.stq_8_bits_succeeded = 1'b1;
    UUT.wrapper.uut.lsu.stq_8_bits_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.lsu.stq_8_bits_uop_dst_rtype = 2'b00;
    UUT.wrapper.uut.lsu.stq_8_bits_uop_exception = 1'b1;
    UUT.wrapper.uut.lsu.stq_8_bits_uop_is_amo = 1'b1;
    UUT.wrapper.uut.lsu.stq_8_bits_uop_is_fence = 1'b1;
    UUT.wrapper.uut.lsu.stq_8_bits_uop_ldq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.stq_8_bits_uop_mem_cmd = 5'b11111;
    UUT.wrapper.uut.lsu.stq_8_bits_uop_mem_signed = 1'b0;
    UUT.wrapper.uut.lsu.stq_8_bits_uop_mem_size = 2'b10;
    UUT.wrapper.uut.lsu.stq_8_bits_uop_pdst = 7'b1111111;
    UUT.wrapper.uut.lsu.stq_8_bits_uop_rob_idx = 6'b000001;
    UUT.wrapper.uut.lsu.stq_8_bits_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.stq_8_bits_uop_uses_ldq = 1'b0;
    UUT.wrapper.uut.lsu.stq_8_bits_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.lsu.stq_8_valid = 1'b1;
    UUT.wrapper.uut.lsu.stq_9_bits_addr_bits = 40'b0000000011111111111111111111100100010111;
    UUT.wrapper.uut.lsu.stq_9_bits_addr_is_virtual = 1'b1;
    UUT.wrapper.uut.lsu.stq_9_bits_addr_valid = 1'b0;
    UUT.wrapper.uut.lsu.stq_9_bits_committed = 1'b1;
    UUT.wrapper.uut.lsu.stq_9_bits_data_bits = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.lsu.stq_9_bits_data_valid = 1'b1;
    UUT.wrapper.uut.lsu.stq_9_bits_debug_wb_data = 64'b1111111111111111111111111111111111111111111111111111111111111111;
    UUT.wrapper.uut.lsu.stq_9_bits_succeeded = 1'b1;
    UUT.wrapper.uut.lsu.stq_9_bits_uop_br_mask = 12'b000000000000;
    UUT.wrapper.uut.lsu.stq_9_bits_uop_dst_rtype = 2'b11;
    UUT.wrapper.uut.lsu.stq_9_bits_uop_exception = 1'b1;
    UUT.wrapper.uut.lsu.stq_9_bits_uop_is_amo = 1'b1;
    UUT.wrapper.uut.lsu.stq_9_bits_uop_is_fence = 1'b1;
    UUT.wrapper.uut.lsu.stq_9_bits_uop_ldq_idx = 4'b1111;
    UUT.wrapper.uut.lsu.stq_9_bits_uop_mem_cmd = 5'b00000;
    UUT.wrapper.uut.lsu.stq_9_bits_uop_mem_signed = 1'b0;
    UUT.wrapper.uut.lsu.stq_9_bits_uop_mem_size = 2'b00;
    UUT.wrapper.uut.lsu.stq_9_bits_uop_pdst = 7'b0000000;
    UUT.wrapper.uut.lsu.stq_9_bits_uop_rob_idx = 6'b111111;
    UUT.wrapper.uut.lsu.stq_9_bits_uop_stq_idx = 4'b0000;
    UUT.wrapper.uut.lsu.stq_9_bits_uop_uses_ldq = 1'b0;
    UUT.wrapper.uut.lsu.stq_9_bits_uop_uses_stq = 1'b0;
    UUT.wrapper.uut.lsu.stq_9_valid = 1'b1;
    UUT.wrapper.uut.lsu.stq_commit_head = 4'b0100;
    UUT.wrapper.uut.lsu.stq_execute_head = 4'b1111;
    UUT.wrapper.uut.lsu.stq_head = 4'b0000;
    UUT.wrapper.uut.lsu.stq_retry_idx = 4'b1111;
    UUT.wrapper.uut.lsu.stq_tail = 4'b0000;
    UUT.wrapper.uut.lsu.wb_forward_ld_addr_0 = 40'b0000000000000000000000000000000000000111;
    UUT.wrapper.uut.lsu.wb_forward_ldq_idx_0 = 4'b1111;
    UUT.wrapper.uut.lsu.wb_forward_stq_idx_0 = 4'b1111;
    UUT.wrapper.uut.lsu.wb_forward_valid_0 = 1'b1;
    UUT.wrapper.uut.ptw.count = 2'b01;
    UUT.wrapper.uut.ptw.l2_refill = 1'b0;
    UUT.wrapper.uut.ptw.mem_resp_data = 64'b0000000000000000000000000000000000000000000000000000001100100001;
    UUT.wrapper.uut.ptw.mem_resp_valid = 1'b1;
    UUT.wrapper.uut.ptw.r_pte_a = 1'b1;
    UUT.wrapper.uut.ptw.r_pte_d = 1'b1;
    UUT.wrapper.uut.ptw.r_pte_g = 1'b1;
    UUT.wrapper.uut.ptw.r_pte_ppn = 44'b11111111111111111111111111111111111111111111;
    UUT.wrapper.uut.ptw.r_pte_r = 1'b1;
    UUT.wrapper.uut.ptw.r_pte_u = 1'b1;
    UUT.wrapper.uut.ptw.r_pte_v = 1'b1;
    UUT.wrapper.uut.ptw.r_pte_w = 1'b1;
    UUT.wrapper.uut.ptw.r_pte_x = 1'b1;
    UUT.wrapper.uut.ptw.r_req_addr = 27'b011111111111110000000001100;
    UUT.wrapper.uut.ptw.r_req_dest = 2'b01;
    UUT.wrapper.uut.ptw.r_req_need_gpa = 1'b0;
    UUT.wrapper.uut.ptw.resp_ae_final = 1'b1;
    UUT.wrapper.uut.ptw.resp_ae_ptw = 1'b1;
    UUT.wrapper.uut.ptw.resp_pf = 1'b1;
    UUT.wrapper.uut.ptw.resp_valid_0 = 1'b1;
    UUT.wrapper.uut.ptw.resp_valid_1 = 1'b1;
    UUT.wrapper.uut.ptw.state = 3'b111;
    UUT.wrapper.uut.tlMasterXbar.beatsLeft = 3'b111;
    UUT.wrapper.uut.tlMasterXbar.readys_mask = 2'b11;
    UUT.wrapper.uut.tlMasterXbar.state_0 = 1'b1;
    UUT.wrapper.uut.tlMasterXbar.state_1 = 1'b1;
    UUT.wrapper.uut.core.rob.rob_debug_wdata[5'b00011] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_debug_wdata[5'b00000] = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    UUT.wrapper.uut.core.rob.rob_debug_wdata[5'b00001] = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    UUT.wrapper.uut.core.rob.rob_debug_wdata[5'b00010] = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    UUT.wrapper.uut.core.rob.rob_debug_wdata_1[5'b00011] = 64'b1000000000000000000000000000000001111111111111111111000000000000;
    UUT.wrapper.uut.core.rob.rob_debug_wdata_1[5'b00000] = 64'b1000000000000000000000000000000001111111111111111111000000000000;
    UUT.wrapper.uut.core.rob.rob_debug_wdata_1[5'b00001] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.core.rob.rob_debug_wdata_1[5'b00010] = 64'b0100000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.dcache.data.array_0_0_0[4'b1110] = 64'b0000000010000000100000000000000001100000000000010000000000000000;
    UUT.wrapper.uut.dcache.meta_0.tag_array_0[1'b1] = 27'b111111111111111110111111111;
    UUT.wrapper.uut.dcache.mshrs.lb[4'b1000] = 64'b0000000000000000000000000000000100000001000000010000000100000001;
    UUT.wrapper.uut.dcache.mshrs.mshrs_0.rpq.ram_addr[1'b1] = 40'b1111111111111111111111111111111111000101;
    UUT.wrapper.uut.dcache.mshrs.mshrs_0.rpq.ram_addr[1'b0] = 40'b0000000000000000000000000000000000111111;
    UUT.wrapper.uut.dcache.mshrs.mshrs_0.rpq.ram_is_hella[1'b1] = 1'b0;
    UUT.wrapper.uut.dcache.mshrs.mshrs_0.rpq.ram_is_hella[1'b0] = 1'b0;
    UUT.wrapper.uut.dcache.mshrs.mshrs_0.rpq.ram_sdq_id[1'b1] = 1'b0;
    UUT.wrapper.uut.dcache.mshrs.mshrs_0.rpq.ram_sdq_id[1'b0] = 1'b1;
    UUT.wrapper.uut.dcache.mshrs.mshrs_1.rpq.ram_addr[1'b1] = 40'b1111111111111111111111111111111110111111;
    UUT.wrapper.uut.dcache.mshrs.mshrs_1.rpq.ram_addr[1'b0] = 40'b1111111111111111111111111111111111101000;
    UUT.wrapper.uut.dcache.mshrs.mshrs_1.rpq.ram_is_hella[1'b1] = 1'b0;
    UUT.wrapper.uut.dcache.mshrs.mshrs_1.rpq.ram_is_hella[1'b0] = 1'b0;
    UUT.wrapper.uut.dcache.mshrs.mshrs_1.rpq.ram_sdq_id[1'b1] = 1'b1;
    UUT.wrapper.uut.dcache.mshrs.mshrs_1.rpq.ram_sdq_id[1'b0] = 1'b1;
    UUT.wrapper.uut.dcache.mshrs.respq.ram_data[2'b11] = 64'b0000000000000000000000000000000000000000000000000000000010100000;
    UUT.wrapper.uut.dcache.mshrs.respq.ram_data[2'b00] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    UUT.wrapper.uut.dcache.mshrs.respq.ram_is_hella[2'b11] = 1'b1;
    UUT.wrapper.uut.dcache.mshrs.respq.ram_is_hella[2'b00] = 1'b0;
    UUT.wrapper.uut.dcache.mshrs.sdq[1'b1] = 64'b0100000010000000100000000000000001010000000000001000000000000000;
    UUT.wrapper.uut.frontend.f3.ram_data[1'b0] = 64'b1001100011000101100111101000001001010111100111011001000001111010;
    UUT.wrapper.uut.frontend.f3.ram_ghist_current_saw_branch_not_taken[1'b0] = 1'b0;
    UUT.wrapper.uut.frontend.f3.ram_ghist_new_saw_branch_not_taken[1'b0] = 1'b0;
    UUT.wrapper.uut.frontend.f3.ram_ghist_new_saw_branch_taken[1'b0] = 1'b1;
    UUT.wrapper.uut.frontend.f3.ram_ghist_old_history[1'b0] = 64'b1110011001100110011001100110011001100110011001100110011001100101;
    UUT.wrapper.uut.frontend.f3.ram_mask[1'b0] = 4'b1010;
    UUT.wrapper.uut.frontend.f3.ram_pc[1'b0] = 40'b0011111111011101110111111111111111111111;
    UUT.wrapper.uut.frontend.f3.ram_xcpt_ae_inst[1'b0] = 1'b1;
    UUT.wrapper.uut.frontend.f3.ram_xcpt_pf_inst[1'b0] = 1'b1;
    UUT.wrapper.uut.frontend.f3_bpd_resp.ram_preds_0_predicted_pc_bits[1'b0] = 40'b0100011101010001110111111111111110110000;
    UUT.wrapper.uut.frontend.f3_bpd_resp.ram_preds_1_predicted_pc_bits[1'b0] = 40'b1111111111111111111111111111111111111111;
    UUT.wrapper.uut.frontend.f3_bpd_resp.ram_preds_2_predicted_pc_bits[1'b0] = 40'b1111111111111111111111111111111111111111;
    UUT.wrapper.uut.frontend.f3_bpd_resp.ram_preds_3_predicted_pc_bits[1'b0] = 40'b1111111111111111111111111111111111111111;
    UUT.wrapper.uut.frontend.f4.ram_bp_debug_if_oh_0[1'b0] = 1'b0;
    UUT.wrapper.uut.frontend.f4.ram_bp_debug_if_oh_1[1'b0] = 1'b0;
    UUT.wrapper.uut.frontend.f4.ram_bp_debug_if_oh_2[1'b0] = 1'b0;
    UUT.wrapper.uut.frontend.f4.ram_bp_debug_if_oh_3[1'b0] = 1'b0;
    UUT.wrapper.uut.frontend.f4.ram_bp_xcpt_if_oh_0[1'b0] = 1'b0;
    UUT.wrapper.uut.frontend.f4.ram_bp_xcpt_if_oh_1[1'b0] = 1'b0;
    UUT.wrapper.uut.frontend.f4.ram_bp_xcpt_if_oh_2[1'b0] = 1'b0;
    UUT.wrapper.uut.frontend.f4.ram_bp_xcpt_if_oh_3[1'b0] = 1'b0;
    UUT.wrapper.uut.frontend.f4.ram_br_mask[1'b0] = 4'b1111;
    UUT.wrapper.uut.frontend.f4.ram_cfi_idx_bits[1'b0] = 2'b11;
    UUT.wrapper.uut.frontend.f4.ram_cfi_idx_valid[1'b0] = 1'b1;
    UUT.wrapper.uut.frontend.f4.ram_edge_inst_0[1'b0] = 1'b0;
    UUT.wrapper.uut.frontend.f4.ram_exp_insts_0[1'b0] = 32'b00000000101001010000001000110011;
    UUT.wrapper.uut.frontend.f4.ram_exp_insts_1[1'b0] = 32'b00000010110000010001010100010011;
    UUT.wrapper.uut.frontend.f4.ram_exp_insts_2[1'b0] = 32'b00111100000001000010001010100011;
    UUT.wrapper.uut.frontend.f4.ram_exp_insts_3[1'b0] = 32'b00000000000000000111000000101011;
    UUT.wrapper.uut.frontend.f4.ram_ghist_current_saw_branch_not_taken[1'b0] = 1'b0;
    UUT.wrapper.uut.frontend.f4.ram_ghist_new_saw_branch_not_taken[1'b0] = 1'b0;
    UUT.wrapper.uut.frontend.f4.ram_ghist_new_saw_branch_taken[1'b0] = 1'b1;
    UUT.wrapper.uut.frontend.f4.ram_ghist_old_history[1'b0] = 64'b1111111111111111111000000001110111011001100110011001100110011000;
    UUT.wrapper.uut.frontend.f4.ram_insts_0[1'b0] = 32'b01000000101001010000011000110111;
    UUT.wrapper.uut.frontend.f4.ram_insts_1[1'b0] = 32'b00100000000010100001000000110010;
    UUT.wrapper.uut.frontend.f4.ram_insts_2[1'b0] = 32'b11000001000000010010001010001110;
    UUT.wrapper.uut.frontend.f4.ram_insts_3[1'b0] = 32'b00000000000000001000000100100011;
    UUT.wrapper.uut.frontend.f4.ram_mask[1'b0] = 4'b1111;
    UUT.wrapper.uut.frontend.f4.ram_pc[1'b0] = 40'b1111100111111010111100111111111111111111;
    UUT.wrapper.uut.frontend.f4.ram_sfbs_0[1'b0] = 1'b1;
    UUT.wrapper.uut.frontend.f4.ram_sfbs_1[1'b0] = 1'b1;
    UUT.wrapper.uut.frontend.f4.ram_sfbs_2[1'b0] = 1'b1;
    UUT.wrapper.uut.frontend.f4.ram_sfbs_3[1'b0] = 1'b0;
    UUT.wrapper.uut.frontend.f4.ram_shadowed_mask_0[1'b0] = 1'b0;
    UUT.wrapper.uut.frontend.f4.ram_shadowed_mask_1[1'b0] = 1'b0;
    UUT.wrapper.uut.frontend.f4.ram_shadowed_mask_2[1'b0] = 1'b0;
    UUT.wrapper.uut.frontend.f4.ram_shadowed_mask_3[1'b0] = 1'b0;
    UUT.wrapper.uut.frontend.f4.ram_xcpt_ae_if[1'b0] = 1'b1;
    UUT.wrapper.uut.frontend.f4.ram_xcpt_pf_if[1'b0] = 1'b0;
    UUT.wrapper.uut.frontend.ftq.ghist_0_current_saw_branch_not_taken[3'b000] = 1'b0;
    UUT.wrapper.uut.frontend.ftq.ghist_0_current_saw_branch_not_taken[3'b010] = 1'b0;
    UUT.wrapper.uut.frontend.ftq.ghist_0_current_saw_branch_not_taken[3'b001] = 1'b0;
    UUT.wrapper.uut.frontend.ftq.ghist_0_old_history[3'b000] = 64'b1011111111111111100000001110111011001100110011001100110011000100;
    UUT.wrapper.uut.frontend.ftq.ghist_0_old_history[3'b010] = 64'b1000111111111111111000000011001100110011001100110011001100110011;
    UUT.wrapper.uut.frontend.ftq.ghist_0_old_history[3'b001] = 64'b0001111111111111110000000110011001100110011001100110011001100110;
    UUT.wrapper.uut.frontend.ftq.ghist_1_current_saw_branch_not_taken[3'b000] = 1'b1;
    UUT.wrapper.uut.frontend.ftq.ghist_1_current_saw_branch_not_taken[3'b001] = 1'b0;
    UUT.wrapper.uut.frontend.ftq.ghist_1_current_saw_branch_not_taken[3'b010] = 1'b0;
    UUT.wrapper.uut.frontend.ftq.ghist_1_new_saw_branch_not_taken[3'b000] = 1'b0;
    UUT.wrapper.uut.frontend.ftq.ghist_1_new_saw_branch_not_taken[3'b001] = 1'b0;
    UUT.wrapper.uut.frontend.ftq.ghist_1_new_saw_branch_not_taken[3'b010] = 1'b0;
    UUT.wrapper.uut.frontend.ftq.ghist_1_new_saw_branch_taken[3'b000] = 1'b0;
    UUT.wrapper.uut.frontend.ftq.ghist_1_new_saw_branch_taken[3'b001] = 1'b0;
    UUT.wrapper.uut.frontend.ftq.ghist_1_new_saw_branch_taken[3'b010] = 1'b0;
    UUT.wrapper.uut.frontend.ftq.ghist_1_old_history[3'b000] = 64'b0001111111111111110000000110011001100110011001100110011001100110;
    UUT.wrapper.uut.frontend.ftq.ghist_1_old_history[3'b001] = 64'b0001111111111111110000000110011001100110011001100110011001100110;
    UUT.wrapper.uut.frontend.ftq.ghist_1_old_history[3'b010] = 64'b0011111111111111100000001100110011001100110011001100110011001100;
    UUT.wrapper.uut.frontend.icache.dataArrayWay_0[4'b1011] = 64'b0100111000100010100011110111111100010011011000001111111001101111;
    UUT.wrapper.uut.frontend.icache.dataArrayWay_0[4'b0000] = 64'b0001001010010111111000001011000110000110000000011000110010000001;
    UUT.wrapper.uut.frontend.icache.dataArrayWay_0[4'b0001] = 64'b1001000000000010111000010000001100100001000100111100000000010001;
    UUT.wrapper.uut.frontend.icache.dataArrayWay_0[4'b0011] = 64'b1110001110001001000111000100000101101101011000110000000100010011;
    UUT.wrapper.uut.frontend.icache.dataArrayWay_0[4'b0010] = 64'b0000000110000011010001100110001110011100010000010110000000010001;
    UUT.wrapper.uut.frontend.icache.dataArrayWay_0[4'b0101] = 64'b1000111011101001000111011010001000101101011000110000000100010011;
    UUT.wrapper.uut.frontend.icache.tag_array_0[1'b0] = 25'b1111111111111111111111111;

    // state 0
    PI_reset = 1'b1;
  end
  always @(posedge clock) begin
    // state 1
    if (cycle == 0) begin
      PI_reset <= 1'b0;
    end

    // state 2
    if (cycle == 1) begin
      PI_reset <= 1'b0;
    end

    // state 3
    if (cycle == 2) begin
      PI_reset <= 1'b0;
    end

    // state 4
    if (cycle == 3) begin
      PI_reset <= 1'b0;
    end

    // state 5
    if (cycle == 4) begin
      PI_reset <= 1'b0;
    end

    // state 6
    if (cycle == 5) begin
      PI_reset <= 1'b0;
    end

    // state 7
    if (cycle == 6) begin
      PI_reset <= 1'b0;
    end

    // state 8
    if (cycle == 7) begin
      PI_reset <= 1'b0;
    end

    // state 9
    if (cycle == 8) begin
      PI_reset <= 1'b0;
    end

    // state 10
    if (cycle == 9) begin
      PI_reset <= 1'b0;
    end

    // state 11
    if (cycle == 10) begin
      PI_reset <= 1'b0;
    end

    // state 12
    if (cycle == 11) begin
      PI_reset <= 1'b0;
    end

    // state 13
    if (cycle == 12) begin
      PI_reset <= 1'b0;
    end

    // state 14
    if (cycle == 13) begin
      PI_reset <= 1'b0;
    end

    // state 15
    if (cycle == 14) begin
      PI_reset <= 1'b0;
    end

    // state 16
    if (cycle == 15) begin
      PI_reset <= 1'b0;
    end

    // state 17
    if (cycle == 16) begin
      PI_reset <= 1'b0;
    end

    // state 18
    if (cycle == 17) begin
      PI_reset <= 1'b0;
    end

    // state 19
    if (cycle == 18) begin
      PI_reset <= 1'b0;
    end

    // state 20
    if (cycle == 19) begin
      PI_reset <= 1'b0;
    end

    genclock <= cycle < 20;
    cycle <= cycle + 1;
  end
endmodule
