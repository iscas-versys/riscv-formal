module SRAMTemplate(
  input         clock,
  input         reset,
  output        io_r_req_ready, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input         io_r_req_valid, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [8:0]  io_r_req_bits_setIdx, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output [27:0] io_r_resp_data_0_tag, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output [1:0]  io_r_resp_data_0__type, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output [38:0] io_r_resp_data_0_target, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output [2:0]  io_r_resp_data_0_brIdx, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output        io_r_resp_data_0_valid, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input         io_w_req_valid, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [8:0]  io_w_req_bits_setIdx, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [27:0] io_w_req_bits_data_tag, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [1:0]  io_w_req_bits_data__type, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [38:0] io_w_req_bits_data_target, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [2:0]  io_w_req_bits_data_brIdx // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [95:0] _RAND_0;
  reg [95:0] _RAND_1;
  reg [95:0] _RAND_2;
  reg [95:0] _RAND_3;
  reg [95:0] _RAND_4;
  reg [95:0] _RAND_5;
  reg [95:0] _RAND_6;
  reg [95:0] _RAND_7;
  reg [95:0] _RAND_8;
  reg [95:0] _RAND_9;
  reg [95:0] _RAND_10;
  reg [95:0] _RAND_11;
  reg [95:0] _RAND_12;
  reg [95:0] _RAND_13;
  reg [95:0] _RAND_14;
  reg [95:0] _RAND_15;
  reg [95:0] _RAND_16;
  reg [95:0] _RAND_17;
  reg [95:0] _RAND_18;
  reg [95:0] _RAND_19;
  reg [95:0] _RAND_20;
  reg [95:0] _RAND_21;
  reg [95:0] _RAND_22;
  reg [95:0] _RAND_23;
  reg [95:0] _RAND_24;
  reg [95:0] _RAND_25;
  reg [95:0] _RAND_26;
  reg [95:0] _RAND_27;
  reg [95:0] _RAND_28;
  reg [95:0] _RAND_29;
  reg [95:0] _RAND_30;
  reg [95:0] _RAND_31;
  reg [95:0] _RAND_32;
  reg [95:0] _RAND_33;
  reg [95:0] _RAND_34;
  reg [95:0] _RAND_35;
  reg [95:0] _RAND_36;
  reg [95:0] _RAND_37;
  reg [95:0] _RAND_38;
  reg [95:0] _RAND_39;
  reg [95:0] _RAND_40;
  reg [95:0] _RAND_41;
  reg [95:0] _RAND_42;
  reg [95:0] _RAND_43;
  reg [95:0] _RAND_44;
  reg [95:0] _RAND_45;
  reg [95:0] _RAND_46;
  reg [95:0] _RAND_47;
  reg [95:0] _RAND_48;
  reg [95:0] _RAND_49;
  reg [95:0] _RAND_50;
  reg [95:0] _RAND_51;
  reg [95:0] _RAND_52;
  reg [95:0] _RAND_53;
  reg [95:0] _RAND_54;
  reg [95:0] _RAND_55;
  reg [95:0] _RAND_56;
  reg [95:0] _RAND_57;
  reg [95:0] _RAND_58;
  reg [95:0] _RAND_59;
  reg [95:0] _RAND_60;
  reg [95:0] _RAND_61;
  reg [95:0] _RAND_62;
  reg [95:0] _RAND_63;
  reg [95:0] _RAND_64;
  reg [95:0] _RAND_65;
  reg [95:0] _RAND_66;
  reg [95:0] _RAND_67;
  reg [95:0] _RAND_68;
  reg [95:0] _RAND_69;
  reg [95:0] _RAND_70;
  reg [95:0] _RAND_71;
  reg [95:0] _RAND_72;
  reg [95:0] _RAND_73;
  reg [95:0] _RAND_74;
  reg [95:0] _RAND_75;
  reg [95:0] _RAND_76;
  reg [95:0] _RAND_77;
  reg [95:0] _RAND_78;
  reg [95:0] _RAND_79;
  reg [95:0] _RAND_80;
  reg [95:0] _RAND_81;
  reg [95:0] _RAND_82;
  reg [95:0] _RAND_83;
  reg [95:0] _RAND_84;
  reg [95:0] _RAND_85;
  reg [95:0] _RAND_86;
  reg [95:0] _RAND_87;
  reg [95:0] _RAND_88;
  reg [95:0] _RAND_89;
  reg [95:0] _RAND_90;
  reg [95:0] _RAND_91;
  reg [95:0] _RAND_92;
  reg [95:0] _RAND_93;
  reg [95:0] _RAND_94;
  reg [95:0] _RAND_95;
  reg [95:0] _RAND_96;
  reg [95:0] _RAND_97;
  reg [95:0] _RAND_98;
  reg [95:0] _RAND_99;
  reg [95:0] _RAND_100;
  reg [95:0] _RAND_101;
  reg [95:0] _RAND_102;
  reg [95:0] _RAND_103;
  reg [95:0] _RAND_104;
  reg [95:0] _RAND_105;
  reg [95:0] _RAND_106;
  reg [95:0] _RAND_107;
  reg [95:0] _RAND_108;
  reg [95:0] _RAND_109;
  reg [95:0] _RAND_110;
  reg [95:0] _RAND_111;
  reg [95:0] _RAND_112;
  reg [95:0] _RAND_113;
  reg [95:0] _RAND_114;
  reg [95:0] _RAND_115;
  reg [95:0] _RAND_116;
  reg [95:0] _RAND_117;
  reg [95:0] _RAND_118;
  reg [95:0] _RAND_119;
  reg [95:0] _RAND_120;
  reg [95:0] _RAND_121;
  reg [95:0] _RAND_122;
  reg [95:0] _RAND_123;
  reg [95:0] _RAND_124;
  reg [95:0] _RAND_125;
  reg [95:0] _RAND_126;
  reg [95:0] _RAND_127;
  reg [95:0] _RAND_128;
  reg [95:0] _RAND_129;
  reg [95:0] _RAND_130;
  reg [95:0] _RAND_131;
  reg [95:0] _RAND_132;
  reg [95:0] _RAND_133;
  reg [95:0] _RAND_134;
  reg [95:0] _RAND_135;
  reg [95:0] _RAND_136;
  reg [95:0] _RAND_137;
  reg [95:0] _RAND_138;
  reg [95:0] _RAND_139;
  reg [95:0] _RAND_140;
  reg [95:0] _RAND_141;
  reg [95:0] _RAND_142;
  reg [95:0] _RAND_143;
  reg [95:0] _RAND_144;
  reg [95:0] _RAND_145;
  reg [95:0] _RAND_146;
  reg [95:0] _RAND_147;
  reg [95:0] _RAND_148;
  reg [95:0] _RAND_149;
  reg [95:0] _RAND_150;
  reg [95:0] _RAND_151;
  reg [95:0] _RAND_152;
  reg [95:0] _RAND_153;
  reg [95:0] _RAND_154;
  reg [95:0] _RAND_155;
  reg [95:0] _RAND_156;
  reg [95:0] _RAND_157;
  reg [95:0] _RAND_158;
  reg [95:0] _RAND_159;
  reg [95:0] _RAND_160;
  reg [95:0] _RAND_161;
  reg [95:0] _RAND_162;
  reg [95:0] _RAND_163;
  reg [95:0] _RAND_164;
  reg [95:0] _RAND_165;
  reg [95:0] _RAND_166;
  reg [95:0] _RAND_167;
  reg [95:0] _RAND_168;
  reg [95:0] _RAND_169;
  reg [95:0] _RAND_170;
  reg [95:0] _RAND_171;
  reg [95:0] _RAND_172;
  reg [95:0] _RAND_173;
  reg [95:0] _RAND_174;
  reg [95:0] _RAND_175;
  reg [95:0] _RAND_176;
  reg [95:0] _RAND_177;
  reg [95:0] _RAND_178;
  reg [95:0] _RAND_179;
  reg [95:0] _RAND_180;
  reg [95:0] _RAND_181;
  reg [95:0] _RAND_182;
  reg [95:0] _RAND_183;
  reg [95:0] _RAND_184;
  reg [95:0] _RAND_185;
  reg [95:0] _RAND_186;
  reg [95:0] _RAND_187;
  reg [95:0] _RAND_188;
  reg [95:0] _RAND_189;
  reg [95:0] _RAND_190;
  reg [95:0] _RAND_191;
  reg [95:0] _RAND_192;
  reg [95:0] _RAND_193;
  reg [95:0] _RAND_194;
  reg [95:0] _RAND_195;
  reg [95:0] _RAND_196;
  reg [95:0] _RAND_197;
  reg [95:0] _RAND_198;
  reg [95:0] _RAND_199;
  reg [95:0] _RAND_200;
  reg [95:0] _RAND_201;
  reg [95:0] _RAND_202;
  reg [95:0] _RAND_203;
  reg [95:0] _RAND_204;
  reg [95:0] _RAND_205;
  reg [95:0] _RAND_206;
  reg [95:0] _RAND_207;
  reg [95:0] _RAND_208;
  reg [95:0] _RAND_209;
  reg [95:0] _RAND_210;
  reg [95:0] _RAND_211;
  reg [95:0] _RAND_212;
  reg [95:0] _RAND_213;
  reg [95:0] _RAND_214;
  reg [95:0] _RAND_215;
  reg [95:0] _RAND_216;
  reg [95:0] _RAND_217;
  reg [95:0] _RAND_218;
  reg [95:0] _RAND_219;
  reg [95:0] _RAND_220;
  reg [95:0] _RAND_221;
  reg [95:0] _RAND_222;
  reg [95:0] _RAND_223;
  reg [95:0] _RAND_224;
  reg [95:0] _RAND_225;
  reg [95:0] _RAND_226;
  reg [95:0] _RAND_227;
  reg [95:0] _RAND_228;
  reg [95:0] _RAND_229;
  reg [95:0] _RAND_230;
  reg [95:0] _RAND_231;
  reg [95:0] _RAND_232;
  reg [95:0] _RAND_233;
  reg [95:0] _RAND_234;
  reg [95:0] _RAND_235;
  reg [95:0] _RAND_236;
  reg [95:0] _RAND_237;
  reg [95:0] _RAND_238;
  reg [95:0] _RAND_239;
  reg [95:0] _RAND_240;
  reg [95:0] _RAND_241;
  reg [95:0] _RAND_242;
  reg [95:0] _RAND_243;
  reg [95:0] _RAND_244;
  reg [95:0] _RAND_245;
  reg [95:0] _RAND_246;
  reg [95:0] _RAND_247;
  reg [95:0] _RAND_248;
  reg [95:0] _RAND_249;
  reg [95:0] _RAND_250;
  reg [95:0] _RAND_251;
  reg [95:0] _RAND_252;
  reg [95:0] _RAND_253;
  reg [95:0] _RAND_254;
  reg [95:0] _RAND_255;
  reg [95:0] _RAND_256;
  reg [95:0] _RAND_257;
  reg [95:0] _RAND_258;
  reg [95:0] _RAND_259;
  reg [95:0] _RAND_260;
  reg [95:0] _RAND_261;
  reg [95:0] _RAND_262;
  reg [95:0] _RAND_263;
  reg [95:0] _RAND_264;
  reg [95:0] _RAND_265;
  reg [95:0] _RAND_266;
  reg [95:0] _RAND_267;
  reg [95:0] _RAND_268;
  reg [95:0] _RAND_269;
  reg [95:0] _RAND_270;
  reg [95:0] _RAND_271;
  reg [95:0] _RAND_272;
  reg [95:0] _RAND_273;
  reg [95:0] _RAND_274;
  reg [95:0] _RAND_275;
  reg [95:0] _RAND_276;
  reg [95:0] _RAND_277;
  reg [95:0] _RAND_278;
  reg [95:0] _RAND_279;
  reg [95:0] _RAND_280;
  reg [95:0] _RAND_281;
  reg [95:0] _RAND_282;
  reg [95:0] _RAND_283;
  reg [95:0] _RAND_284;
  reg [95:0] _RAND_285;
  reg [95:0] _RAND_286;
  reg [95:0] _RAND_287;
  reg [95:0] _RAND_288;
  reg [95:0] _RAND_289;
  reg [95:0] _RAND_290;
  reg [95:0] _RAND_291;
  reg [95:0] _RAND_292;
  reg [95:0] _RAND_293;
  reg [95:0] _RAND_294;
  reg [95:0] _RAND_295;
  reg [95:0] _RAND_296;
  reg [95:0] _RAND_297;
  reg [95:0] _RAND_298;
  reg [95:0] _RAND_299;
  reg [95:0] _RAND_300;
  reg [95:0] _RAND_301;
  reg [95:0] _RAND_302;
  reg [95:0] _RAND_303;
  reg [95:0] _RAND_304;
  reg [95:0] _RAND_305;
  reg [95:0] _RAND_306;
  reg [95:0] _RAND_307;
  reg [95:0] _RAND_308;
  reg [95:0] _RAND_309;
  reg [95:0] _RAND_310;
  reg [95:0] _RAND_311;
  reg [95:0] _RAND_312;
  reg [95:0] _RAND_313;
  reg [95:0] _RAND_314;
  reg [95:0] _RAND_315;
  reg [95:0] _RAND_316;
  reg [95:0] _RAND_317;
  reg [95:0] _RAND_318;
  reg [95:0] _RAND_319;
  reg [95:0] _RAND_320;
  reg [95:0] _RAND_321;
  reg [95:0] _RAND_322;
  reg [95:0] _RAND_323;
  reg [95:0] _RAND_324;
  reg [95:0] _RAND_325;
  reg [95:0] _RAND_326;
  reg [95:0] _RAND_327;
  reg [95:0] _RAND_328;
  reg [95:0] _RAND_329;
  reg [95:0] _RAND_330;
  reg [95:0] _RAND_331;
  reg [95:0] _RAND_332;
  reg [95:0] _RAND_333;
  reg [95:0] _RAND_334;
  reg [95:0] _RAND_335;
  reg [95:0] _RAND_336;
  reg [95:0] _RAND_337;
  reg [95:0] _RAND_338;
  reg [95:0] _RAND_339;
  reg [95:0] _RAND_340;
  reg [95:0] _RAND_341;
  reg [95:0] _RAND_342;
  reg [95:0] _RAND_343;
  reg [95:0] _RAND_344;
  reg [95:0] _RAND_345;
  reg [95:0] _RAND_346;
  reg [95:0] _RAND_347;
  reg [95:0] _RAND_348;
  reg [95:0] _RAND_349;
  reg [95:0] _RAND_350;
  reg [95:0] _RAND_351;
  reg [95:0] _RAND_352;
  reg [95:0] _RAND_353;
  reg [95:0] _RAND_354;
  reg [95:0] _RAND_355;
  reg [95:0] _RAND_356;
  reg [95:0] _RAND_357;
  reg [95:0] _RAND_358;
  reg [95:0] _RAND_359;
  reg [95:0] _RAND_360;
  reg [95:0] _RAND_361;
  reg [95:0] _RAND_362;
  reg [95:0] _RAND_363;
  reg [95:0] _RAND_364;
  reg [95:0] _RAND_365;
  reg [95:0] _RAND_366;
  reg [95:0] _RAND_367;
  reg [95:0] _RAND_368;
  reg [95:0] _RAND_369;
  reg [95:0] _RAND_370;
  reg [95:0] _RAND_371;
  reg [95:0] _RAND_372;
  reg [95:0] _RAND_373;
  reg [95:0] _RAND_374;
  reg [95:0] _RAND_375;
  reg [95:0] _RAND_376;
  reg [95:0] _RAND_377;
  reg [95:0] _RAND_378;
  reg [95:0] _RAND_379;
  reg [95:0] _RAND_380;
  reg [95:0] _RAND_381;
  reg [95:0] _RAND_382;
  reg [95:0] _RAND_383;
  reg [95:0] _RAND_384;
  reg [95:0] _RAND_385;
  reg [95:0] _RAND_386;
  reg [95:0] _RAND_387;
  reg [95:0] _RAND_388;
  reg [95:0] _RAND_389;
  reg [95:0] _RAND_390;
  reg [95:0] _RAND_391;
  reg [95:0] _RAND_392;
  reg [95:0] _RAND_393;
  reg [95:0] _RAND_394;
  reg [95:0] _RAND_395;
  reg [95:0] _RAND_396;
  reg [95:0] _RAND_397;
  reg [95:0] _RAND_398;
  reg [95:0] _RAND_399;
  reg [95:0] _RAND_400;
  reg [95:0] _RAND_401;
  reg [95:0] _RAND_402;
  reg [95:0] _RAND_403;
  reg [95:0] _RAND_404;
  reg [95:0] _RAND_405;
  reg [95:0] _RAND_406;
  reg [95:0] _RAND_407;
  reg [95:0] _RAND_408;
  reg [95:0] _RAND_409;
  reg [95:0] _RAND_410;
  reg [95:0] _RAND_411;
  reg [95:0] _RAND_412;
  reg [95:0] _RAND_413;
  reg [95:0] _RAND_414;
  reg [95:0] _RAND_415;
  reg [95:0] _RAND_416;
  reg [95:0] _RAND_417;
  reg [95:0] _RAND_418;
  reg [95:0] _RAND_419;
  reg [95:0] _RAND_420;
  reg [95:0] _RAND_421;
  reg [95:0] _RAND_422;
  reg [95:0] _RAND_423;
  reg [95:0] _RAND_424;
  reg [95:0] _RAND_425;
  reg [95:0] _RAND_426;
  reg [95:0] _RAND_427;
  reg [95:0] _RAND_428;
  reg [95:0] _RAND_429;
  reg [95:0] _RAND_430;
  reg [95:0] _RAND_431;
  reg [95:0] _RAND_432;
  reg [95:0] _RAND_433;
  reg [95:0] _RAND_434;
  reg [95:0] _RAND_435;
  reg [95:0] _RAND_436;
  reg [95:0] _RAND_437;
  reg [95:0] _RAND_438;
  reg [95:0] _RAND_439;
  reg [95:0] _RAND_440;
  reg [95:0] _RAND_441;
  reg [95:0] _RAND_442;
  reg [95:0] _RAND_443;
  reg [95:0] _RAND_444;
  reg [95:0] _RAND_445;
  reg [95:0] _RAND_446;
  reg [95:0] _RAND_447;
  reg [95:0] _RAND_448;
  reg [95:0] _RAND_449;
  reg [95:0] _RAND_450;
  reg [95:0] _RAND_451;
  reg [95:0] _RAND_452;
  reg [95:0] _RAND_453;
  reg [95:0] _RAND_454;
  reg [95:0] _RAND_455;
  reg [95:0] _RAND_456;
  reg [95:0] _RAND_457;
  reg [95:0] _RAND_458;
  reg [95:0] _RAND_459;
  reg [95:0] _RAND_460;
  reg [95:0] _RAND_461;
  reg [95:0] _RAND_462;
  reg [95:0] _RAND_463;
  reg [95:0] _RAND_464;
  reg [95:0] _RAND_465;
  reg [95:0] _RAND_466;
  reg [95:0] _RAND_467;
  reg [95:0] _RAND_468;
  reg [95:0] _RAND_469;
  reg [95:0] _RAND_470;
  reg [95:0] _RAND_471;
  reg [95:0] _RAND_472;
  reg [95:0] _RAND_473;
  reg [95:0] _RAND_474;
  reg [95:0] _RAND_475;
  reg [95:0] _RAND_476;
  reg [95:0] _RAND_477;
  reg [95:0] _RAND_478;
  reg [95:0] _RAND_479;
  reg [95:0] _RAND_480;
  reg [95:0] _RAND_481;
  reg [95:0] _RAND_482;
  reg [95:0] _RAND_483;
  reg [95:0] _RAND_484;
  reg [95:0] _RAND_485;
  reg [95:0] _RAND_486;
  reg [95:0] _RAND_487;
  reg [95:0] _RAND_488;
  reg [95:0] _RAND_489;
  reg [95:0] _RAND_490;
  reg [95:0] _RAND_491;
  reg [95:0] _RAND_492;
  reg [95:0] _RAND_493;
  reg [95:0] _RAND_494;
  reg [95:0] _RAND_495;
  reg [95:0] _RAND_496;
  reg [95:0] _RAND_497;
  reg [95:0] _RAND_498;
  reg [95:0] _RAND_499;
  reg [95:0] _RAND_500;
  reg [95:0] _RAND_501;
  reg [95:0] _RAND_502;
  reg [95:0] _RAND_503;
  reg [95:0] _RAND_504;
  reg [95:0] _RAND_505;
  reg [95:0] _RAND_506;
  reg [95:0] _RAND_507;
  reg [95:0] _RAND_508;
  reg [95:0] _RAND_509;
  reg [95:0] _RAND_510;
  reg [95:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [95:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [95:0] _RAND_516;
`endif // RANDOMIZE_REG_INIT
  reg [72:0] regs_0_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_1_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_2_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_3_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_4_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_5_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_6_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_7_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_8_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_9_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_10_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_11_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_12_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_13_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_14_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_15_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_16_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_17_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_18_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_19_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_20_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_21_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_22_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_23_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_24_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_25_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_26_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_27_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_28_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_29_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_30_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_31_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_32_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_33_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_34_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_35_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_36_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_37_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_38_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_39_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_40_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_41_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_42_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_43_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_44_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_45_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_46_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_47_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_48_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_49_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_50_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_51_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_52_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_53_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_54_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_55_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_56_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_57_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_58_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_59_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_60_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_61_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_62_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_63_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_64_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_65_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_66_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_67_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_68_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_69_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_70_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_71_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_72_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_73_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_74_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_75_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_76_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_77_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_78_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_79_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_80_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_81_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_82_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_83_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_84_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_85_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_86_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_87_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_88_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_89_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_90_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_91_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_92_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_93_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_94_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_95_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_96_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_97_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_98_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_99_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_100_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_101_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_102_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_103_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_104_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_105_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_106_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_107_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_108_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_109_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_110_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_111_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_112_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_113_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_114_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_115_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_116_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_117_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_118_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_119_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_120_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_121_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_122_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_123_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_124_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_125_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_126_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_127_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_128_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_129_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_130_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_131_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_132_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_133_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_134_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_135_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_136_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_137_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_138_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_139_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_140_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_141_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_142_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_143_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_144_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_145_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_146_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_147_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_148_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_149_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_150_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_151_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_152_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_153_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_154_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_155_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_156_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_157_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_158_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_159_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_160_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_161_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_162_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_163_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_164_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_165_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_166_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_167_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_168_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_169_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_170_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_171_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_172_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_173_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_174_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_175_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_176_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_177_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_178_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_179_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_180_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_181_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_182_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_183_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_184_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_185_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_186_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_187_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_188_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_189_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_190_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_191_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_192_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_193_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_194_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_195_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_196_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_197_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_198_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_199_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_200_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_201_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_202_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_203_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_204_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_205_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_206_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_207_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_208_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_209_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_210_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_211_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_212_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_213_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_214_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_215_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_216_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_217_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_218_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_219_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_220_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_221_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_222_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_223_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_224_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_225_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_226_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_227_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_228_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_229_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_230_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_231_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_232_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_233_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_234_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_235_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_236_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_237_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_238_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_239_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_240_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_241_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_242_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_243_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_244_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_245_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_246_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_247_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_248_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_249_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_250_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_251_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_252_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_253_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_254_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_255_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_256_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_257_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_258_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_259_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_260_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_261_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_262_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_263_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_264_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_265_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_266_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_267_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_268_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_269_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_270_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_271_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_272_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_273_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_274_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_275_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_276_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_277_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_278_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_279_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_280_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_281_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_282_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_283_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_284_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_285_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_286_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_287_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_288_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_289_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_290_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_291_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_292_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_293_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_294_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_295_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_296_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_297_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_298_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_299_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_300_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_301_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_302_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_303_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_304_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_305_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_306_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_307_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_308_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_309_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_310_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_311_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_312_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_313_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_314_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_315_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_316_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_317_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_318_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_319_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_320_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_321_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_322_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_323_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_324_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_325_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_326_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_327_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_328_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_329_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_330_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_331_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_332_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_333_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_334_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_335_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_336_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_337_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_338_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_339_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_340_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_341_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_342_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_343_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_344_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_345_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_346_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_347_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_348_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_349_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_350_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_351_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_352_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_353_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_354_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_355_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_356_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_357_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_358_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_359_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_360_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_361_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_362_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_363_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_364_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_365_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_366_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_367_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_368_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_369_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_370_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_371_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_372_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_373_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_374_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_375_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_376_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_377_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_378_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_379_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_380_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_381_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_382_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_383_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_384_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_385_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_386_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_387_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_388_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_389_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_390_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_391_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_392_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_393_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_394_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_395_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_396_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_397_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_398_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_399_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_400_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_401_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_402_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_403_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_404_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_405_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_406_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_407_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_408_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_409_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_410_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_411_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_412_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_413_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_414_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_415_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_416_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_417_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_418_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_419_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_420_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_421_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_422_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_423_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_424_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_425_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_426_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_427_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_428_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_429_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_430_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_431_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_432_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_433_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_434_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_435_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_436_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_437_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_438_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_439_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_440_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_441_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_442_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_443_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_444_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_445_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_446_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_447_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_448_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_449_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_450_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_451_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_452_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_453_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_454_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_455_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_456_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_457_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_458_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_459_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_460_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_461_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_462_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_463_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_464_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_465_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_466_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_467_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_468_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_469_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_470_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_471_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_472_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_473_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_474_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_475_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_476_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_477_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_478_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_479_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_480_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_481_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_482_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_483_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_484_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_485_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_486_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_487_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_488_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_489_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_490_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_491_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_492_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_493_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_494_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_495_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_496_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_497_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_498_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_499_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_500_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_501_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_502_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_503_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_504_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_505_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_506_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_507_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_508_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_509_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_510_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [72:0] regs_511_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg  resetState; // @[src/main/scala/utils/SRAMTemplate.scala 80:30]
  reg [8:0] resetSet; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  wrap_wrap = resetSet == 9'h1ff; // @[src/main/scala/chisel3/util/Counter.scala 73:24]
  wire [8:0] _wrap_value_T_1 = resetSet + 9'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  resetFinish = resetState & wrap_wrap; // @[src/main/scala/chisel3/util/Counter.scala 118:{16,23} 117:24]
  wire  _GEN_2 = resetFinish ? 1'h0 : resetState; // @[src/main/scala/utils/SRAMTemplate.scala 82:24 80:30 82:38]
  wire  wen = io_w_req_valid | resetState; // @[src/main/scala/utils/SRAMTemplate.scala 88:52]
  wire  _realRen_T = ~wen; // @[src/main/scala/utils/SRAMTemplate.scala 89:41]
  wire  realRen = io_r_req_valid & ~wen; // @[src/main/scala/utils/SRAMTemplate.scala 89:38]
  wire [8:0] setIdx = resetState ? resetSet : io_w_req_bits_setIdx; // @[src/main/scala/utils/SRAMTemplate.scala 91:19]
  wire [72:0] _wdataword_T = {io_w_req_bits_data_tag,io_w_req_bits_data__type,io_w_req_bits_data_target,
    io_w_req_bits_data_brIdx,1'h1}; // @[src/main/scala/utils/SRAMTemplate.scala 92:78]
  reg [72:0] rdata_r_0; // @[src/main/scala/utils/RegMem.scala 39:14]
  wire [72:0] _GEN_1540 = 9'h1 == io_r_req_bits_setIdx ? regs_1_0 : regs_0_0; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1541 = 9'h2 == io_r_req_bits_setIdx ? regs_2_0 : _GEN_1540; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1542 = 9'h3 == io_r_req_bits_setIdx ? regs_3_0 : _GEN_1541; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1543 = 9'h4 == io_r_req_bits_setIdx ? regs_4_0 : _GEN_1542; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1544 = 9'h5 == io_r_req_bits_setIdx ? regs_5_0 : _GEN_1543; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1545 = 9'h6 == io_r_req_bits_setIdx ? regs_6_0 : _GEN_1544; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1546 = 9'h7 == io_r_req_bits_setIdx ? regs_7_0 : _GEN_1545; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1547 = 9'h8 == io_r_req_bits_setIdx ? regs_8_0 : _GEN_1546; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1548 = 9'h9 == io_r_req_bits_setIdx ? regs_9_0 : _GEN_1547; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1549 = 9'ha == io_r_req_bits_setIdx ? regs_10_0 : _GEN_1548; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1550 = 9'hb == io_r_req_bits_setIdx ? regs_11_0 : _GEN_1549; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1551 = 9'hc == io_r_req_bits_setIdx ? regs_12_0 : _GEN_1550; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1552 = 9'hd == io_r_req_bits_setIdx ? regs_13_0 : _GEN_1551; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1553 = 9'he == io_r_req_bits_setIdx ? regs_14_0 : _GEN_1552; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1554 = 9'hf == io_r_req_bits_setIdx ? regs_15_0 : _GEN_1553; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1555 = 9'h10 == io_r_req_bits_setIdx ? regs_16_0 : _GEN_1554; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1556 = 9'h11 == io_r_req_bits_setIdx ? regs_17_0 : _GEN_1555; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1557 = 9'h12 == io_r_req_bits_setIdx ? regs_18_0 : _GEN_1556; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1558 = 9'h13 == io_r_req_bits_setIdx ? regs_19_0 : _GEN_1557; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1559 = 9'h14 == io_r_req_bits_setIdx ? regs_20_0 : _GEN_1558; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1560 = 9'h15 == io_r_req_bits_setIdx ? regs_21_0 : _GEN_1559; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1561 = 9'h16 == io_r_req_bits_setIdx ? regs_22_0 : _GEN_1560; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1562 = 9'h17 == io_r_req_bits_setIdx ? regs_23_0 : _GEN_1561; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1563 = 9'h18 == io_r_req_bits_setIdx ? regs_24_0 : _GEN_1562; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1564 = 9'h19 == io_r_req_bits_setIdx ? regs_25_0 : _GEN_1563; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1565 = 9'h1a == io_r_req_bits_setIdx ? regs_26_0 : _GEN_1564; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1566 = 9'h1b == io_r_req_bits_setIdx ? regs_27_0 : _GEN_1565; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1567 = 9'h1c == io_r_req_bits_setIdx ? regs_28_0 : _GEN_1566; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1568 = 9'h1d == io_r_req_bits_setIdx ? regs_29_0 : _GEN_1567; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1569 = 9'h1e == io_r_req_bits_setIdx ? regs_30_0 : _GEN_1568; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1570 = 9'h1f == io_r_req_bits_setIdx ? regs_31_0 : _GEN_1569; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1571 = 9'h20 == io_r_req_bits_setIdx ? regs_32_0 : _GEN_1570; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1572 = 9'h21 == io_r_req_bits_setIdx ? regs_33_0 : _GEN_1571; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1573 = 9'h22 == io_r_req_bits_setIdx ? regs_34_0 : _GEN_1572; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1574 = 9'h23 == io_r_req_bits_setIdx ? regs_35_0 : _GEN_1573; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1575 = 9'h24 == io_r_req_bits_setIdx ? regs_36_0 : _GEN_1574; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1576 = 9'h25 == io_r_req_bits_setIdx ? regs_37_0 : _GEN_1575; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1577 = 9'h26 == io_r_req_bits_setIdx ? regs_38_0 : _GEN_1576; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1578 = 9'h27 == io_r_req_bits_setIdx ? regs_39_0 : _GEN_1577; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1579 = 9'h28 == io_r_req_bits_setIdx ? regs_40_0 : _GEN_1578; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1580 = 9'h29 == io_r_req_bits_setIdx ? regs_41_0 : _GEN_1579; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1581 = 9'h2a == io_r_req_bits_setIdx ? regs_42_0 : _GEN_1580; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1582 = 9'h2b == io_r_req_bits_setIdx ? regs_43_0 : _GEN_1581; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1583 = 9'h2c == io_r_req_bits_setIdx ? regs_44_0 : _GEN_1582; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1584 = 9'h2d == io_r_req_bits_setIdx ? regs_45_0 : _GEN_1583; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1585 = 9'h2e == io_r_req_bits_setIdx ? regs_46_0 : _GEN_1584; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1586 = 9'h2f == io_r_req_bits_setIdx ? regs_47_0 : _GEN_1585; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1587 = 9'h30 == io_r_req_bits_setIdx ? regs_48_0 : _GEN_1586; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1588 = 9'h31 == io_r_req_bits_setIdx ? regs_49_0 : _GEN_1587; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1589 = 9'h32 == io_r_req_bits_setIdx ? regs_50_0 : _GEN_1588; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1590 = 9'h33 == io_r_req_bits_setIdx ? regs_51_0 : _GEN_1589; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1591 = 9'h34 == io_r_req_bits_setIdx ? regs_52_0 : _GEN_1590; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1592 = 9'h35 == io_r_req_bits_setIdx ? regs_53_0 : _GEN_1591; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1593 = 9'h36 == io_r_req_bits_setIdx ? regs_54_0 : _GEN_1592; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1594 = 9'h37 == io_r_req_bits_setIdx ? regs_55_0 : _GEN_1593; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1595 = 9'h38 == io_r_req_bits_setIdx ? regs_56_0 : _GEN_1594; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1596 = 9'h39 == io_r_req_bits_setIdx ? regs_57_0 : _GEN_1595; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1597 = 9'h3a == io_r_req_bits_setIdx ? regs_58_0 : _GEN_1596; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1598 = 9'h3b == io_r_req_bits_setIdx ? regs_59_0 : _GEN_1597; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1599 = 9'h3c == io_r_req_bits_setIdx ? regs_60_0 : _GEN_1598; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1600 = 9'h3d == io_r_req_bits_setIdx ? regs_61_0 : _GEN_1599; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1601 = 9'h3e == io_r_req_bits_setIdx ? regs_62_0 : _GEN_1600; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1602 = 9'h3f == io_r_req_bits_setIdx ? regs_63_0 : _GEN_1601; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1603 = 9'h40 == io_r_req_bits_setIdx ? regs_64_0 : _GEN_1602; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1604 = 9'h41 == io_r_req_bits_setIdx ? regs_65_0 : _GEN_1603; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1605 = 9'h42 == io_r_req_bits_setIdx ? regs_66_0 : _GEN_1604; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1606 = 9'h43 == io_r_req_bits_setIdx ? regs_67_0 : _GEN_1605; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1607 = 9'h44 == io_r_req_bits_setIdx ? regs_68_0 : _GEN_1606; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1608 = 9'h45 == io_r_req_bits_setIdx ? regs_69_0 : _GEN_1607; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1609 = 9'h46 == io_r_req_bits_setIdx ? regs_70_0 : _GEN_1608; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1610 = 9'h47 == io_r_req_bits_setIdx ? regs_71_0 : _GEN_1609; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1611 = 9'h48 == io_r_req_bits_setIdx ? regs_72_0 : _GEN_1610; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1612 = 9'h49 == io_r_req_bits_setIdx ? regs_73_0 : _GEN_1611; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1613 = 9'h4a == io_r_req_bits_setIdx ? regs_74_0 : _GEN_1612; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1614 = 9'h4b == io_r_req_bits_setIdx ? regs_75_0 : _GEN_1613; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1615 = 9'h4c == io_r_req_bits_setIdx ? regs_76_0 : _GEN_1614; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1616 = 9'h4d == io_r_req_bits_setIdx ? regs_77_0 : _GEN_1615; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1617 = 9'h4e == io_r_req_bits_setIdx ? regs_78_0 : _GEN_1616; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1618 = 9'h4f == io_r_req_bits_setIdx ? regs_79_0 : _GEN_1617; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1619 = 9'h50 == io_r_req_bits_setIdx ? regs_80_0 : _GEN_1618; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1620 = 9'h51 == io_r_req_bits_setIdx ? regs_81_0 : _GEN_1619; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1621 = 9'h52 == io_r_req_bits_setIdx ? regs_82_0 : _GEN_1620; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1622 = 9'h53 == io_r_req_bits_setIdx ? regs_83_0 : _GEN_1621; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1623 = 9'h54 == io_r_req_bits_setIdx ? regs_84_0 : _GEN_1622; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1624 = 9'h55 == io_r_req_bits_setIdx ? regs_85_0 : _GEN_1623; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1625 = 9'h56 == io_r_req_bits_setIdx ? regs_86_0 : _GEN_1624; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1626 = 9'h57 == io_r_req_bits_setIdx ? regs_87_0 : _GEN_1625; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1627 = 9'h58 == io_r_req_bits_setIdx ? regs_88_0 : _GEN_1626; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1628 = 9'h59 == io_r_req_bits_setIdx ? regs_89_0 : _GEN_1627; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1629 = 9'h5a == io_r_req_bits_setIdx ? regs_90_0 : _GEN_1628; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1630 = 9'h5b == io_r_req_bits_setIdx ? regs_91_0 : _GEN_1629; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1631 = 9'h5c == io_r_req_bits_setIdx ? regs_92_0 : _GEN_1630; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1632 = 9'h5d == io_r_req_bits_setIdx ? regs_93_0 : _GEN_1631; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1633 = 9'h5e == io_r_req_bits_setIdx ? regs_94_0 : _GEN_1632; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1634 = 9'h5f == io_r_req_bits_setIdx ? regs_95_0 : _GEN_1633; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1635 = 9'h60 == io_r_req_bits_setIdx ? regs_96_0 : _GEN_1634; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1636 = 9'h61 == io_r_req_bits_setIdx ? regs_97_0 : _GEN_1635; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1637 = 9'h62 == io_r_req_bits_setIdx ? regs_98_0 : _GEN_1636; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1638 = 9'h63 == io_r_req_bits_setIdx ? regs_99_0 : _GEN_1637; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1639 = 9'h64 == io_r_req_bits_setIdx ? regs_100_0 : _GEN_1638; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1640 = 9'h65 == io_r_req_bits_setIdx ? regs_101_0 : _GEN_1639; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1641 = 9'h66 == io_r_req_bits_setIdx ? regs_102_0 : _GEN_1640; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1642 = 9'h67 == io_r_req_bits_setIdx ? regs_103_0 : _GEN_1641; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1643 = 9'h68 == io_r_req_bits_setIdx ? regs_104_0 : _GEN_1642; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1644 = 9'h69 == io_r_req_bits_setIdx ? regs_105_0 : _GEN_1643; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1645 = 9'h6a == io_r_req_bits_setIdx ? regs_106_0 : _GEN_1644; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1646 = 9'h6b == io_r_req_bits_setIdx ? regs_107_0 : _GEN_1645; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1647 = 9'h6c == io_r_req_bits_setIdx ? regs_108_0 : _GEN_1646; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1648 = 9'h6d == io_r_req_bits_setIdx ? regs_109_0 : _GEN_1647; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1649 = 9'h6e == io_r_req_bits_setIdx ? regs_110_0 : _GEN_1648; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1650 = 9'h6f == io_r_req_bits_setIdx ? regs_111_0 : _GEN_1649; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1651 = 9'h70 == io_r_req_bits_setIdx ? regs_112_0 : _GEN_1650; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1652 = 9'h71 == io_r_req_bits_setIdx ? regs_113_0 : _GEN_1651; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1653 = 9'h72 == io_r_req_bits_setIdx ? regs_114_0 : _GEN_1652; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1654 = 9'h73 == io_r_req_bits_setIdx ? regs_115_0 : _GEN_1653; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1655 = 9'h74 == io_r_req_bits_setIdx ? regs_116_0 : _GEN_1654; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1656 = 9'h75 == io_r_req_bits_setIdx ? regs_117_0 : _GEN_1655; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1657 = 9'h76 == io_r_req_bits_setIdx ? regs_118_0 : _GEN_1656; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1658 = 9'h77 == io_r_req_bits_setIdx ? regs_119_0 : _GEN_1657; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1659 = 9'h78 == io_r_req_bits_setIdx ? regs_120_0 : _GEN_1658; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1660 = 9'h79 == io_r_req_bits_setIdx ? regs_121_0 : _GEN_1659; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1661 = 9'h7a == io_r_req_bits_setIdx ? regs_122_0 : _GEN_1660; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1662 = 9'h7b == io_r_req_bits_setIdx ? regs_123_0 : _GEN_1661; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1663 = 9'h7c == io_r_req_bits_setIdx ? regs_124_0 : _GEN_1662; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1664 = 9'h7d == io_r_req_bits_setIdx ? regs_125_0 : _GEN_1663; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1665 = 9'h7e == io_r_req_bits_setIdx ? regs_126_0 : _GEN_1664; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1666 = 9'h7f == io_r_req_bits_setIdx ? regs_127_0 : _GEN_1665; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1667 = 9'h80 == io_r_req_bits_setIdx ? regs_128_0 : _GEN_1666; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1668 = 9'h81 == io_r_req_bits_setIdx ? regs_129_0 : _GEN_1667; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1669 = 9'h82 == io_r_req_bits_setIdx ? regs_130_0 : _GEN_1668; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1670 = 9'h83 == io_r_req_bits_setIdx ? regs_131_0 : _GEN_1669; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1671 = 9'h84 == io_r_req_bits_setIdx ? regs_132_0 : _GEN_1670; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1672 = 9'h85 == io_r_req_bits_setIdx ? regs_133_0 : _GEN_1671; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1673 = 9'h86 == io_r_req_bits_setIdx ? regs_134_0 : _GEN_1672; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1674 = 9'h87 == io_r_req_bits_setIdx ? regs_135_0 : _GEN_1673; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1675 = 9'h88 == io_r_req_bits_setIdx ? regs_136_0 : _GEN_1674; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1676 = 9'h89 == io_r_req_bits_setIdx ? regs_137_0 : _GEN_1675; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1677 = 9'h8a == io_r_req_bits_setIdx ? regs_138_0 : _GEN_1676; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1678 = 9'h8b == io_r_req_bits_setIdx ? regs_139_0 : _GEN_1677; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1679 = 9'h8c == io_r_req_bits_setIdx ? regs_140_0 : _GEN_1678; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1680 = 9'h8d == io_r_req_bits_setIdx ? regs_141_0 : _GEN_1679; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1681 = 9'h8e == io_r_req_bits_setIdx ? regs_142_0 : _GEN_1680; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1682 = 9'h8f == io_r_req_bits_setIdx ? regs_143_0 : _GEN_1681; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1683 = 9'h90 == io_r_req_bits_setIdx ? regs_144_0 : _GEN_1682; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1684 = 9'h91 == io_r_req_bits_setIdx ? regs_145_0 : _GEN_1683; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1685 = 9'h92 == io_r_req_bits_setIdx ? regs_146_0 : _GEN_1684; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1686 = 9'h93 == io_r_req_bits_setIdx ? regs_147_0 : _GEN_1685; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1687 = 9'h94 == io_r_req_bits_setIdx ? regs_148_0 : _GEN_1686; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1688 = 9'h95 == io_r_req_bits_setIdx ? regs_149_0 : _GEN_1687; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1689 = 9'h96 == io_r_req_bits_setIdx ? regs_150_0 : _GEN_1688; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1690 = 9'h97 == io_r_req_bits_setIdx ? regs_151_0 : _GEN_1689; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1691 = 9'h98 == io_r_req_bits_setIdx ? regs_152_0 : _GEN_1690; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1692 = 9'h99 == io_r_req_bits_setIdx ? regs_153_0 : _GEN_1691; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1693 = 9'h9a == io_r_req_bits_setIdx ? regs_154_0 : _GEN_1692; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1694 = 9'h9b == io_r_req_bits_setIdx ? regs_155_0 : _GEN_1693; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1695 = 9'h9c == io_r_req_bits_setIdx ? regs_156_0 : _GEN_1694; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1696 = 9'h9d == io_r_req_bits_setIdx ? regs_157_0 : _GEN_1695; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1697 = 9'h9e == io_r_req_bits_setIdx ? regs_158_0 : _GEN_1696; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1698 = 9'h9f == io_r_req_bits_setIdx ? regs_159_0 : _GEN_1697; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1699 = 9'ha0 == io_r_req_bits_setIdx ? regs_160_0 : _GEN_1698; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1700 = 9'ha1 == io_r_req_bits_setIdx ? regs_161_0 : _GEN_1699; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1701 = 9'ha2 == io_r_req_bits_setIdx ? regs_162_0 : _GEN_1700; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1702 = 9'ha3 == io_r_req_bits_setIdx ? regs_163_0 : _GEN_1701; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1703 = 9'ha4 == io_r_req_bits_setIdx ? regs_164_0 : _GEN_1702; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1704 = 9'ha5 == io_r_req_bits_setIdx ? regs_165_0 : _GEN_1703; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1705 = 9'ha6 == io_r_req_bits_setIdx ? regs_166_0 : _GEN_1704; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1706 = 9'ha7 == io_r_req_bits_setIdx ? regs_167_0 : _GEN_1705; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1707 = 9'ha8 == io_r_req_bits_setIdx ? regs_168_0 : _GEN_1706; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1708 = 9'ha9 == io_r_req_bits_setIdx ? regs_169_0 : _GEN_1707; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1709 = 9'haa == io_r_req_bits_setIdx ? regs_170_0 : _GEN_1708; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1710 = 9'hab == io_r_req_bits_setIdx ? regs_171_0 : _GEN_1709; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1711 = 9'hac == io_r_req_bits_setIdx ? regs_172_0 : _GEN_1710; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1712 = 9'had == io_r_req_bits_setIdx ? regs_173_0 : _GEN_1711; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1713 = 9'hae == io_r_req_bits_setIdx ? regs_174_0 : _GEN_1712; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1714 = 9'haf == io_r_req_bits_setIdx ? regs_175_0 : _GEN_1713; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1715 = 9'hb0 == io_r_req_bits_setIdx ? regs_176_0 : _GEN_1714; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1716 = 9'hb1 == io_r_req_bits_setIdx ? regs_177_0 : _GEN_1715; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1717 = 9'hb2 == io_r_req_bits_setIdx ? regs_178_0 : _GEN_1716; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1718 = 9'hb3 == io_r_req_bits_setIdx ? regs_179_0 : _GEN_1717; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1719 = 9'hb4 == io_r_req_bits_setIdx ? regs_180_0 : _GEN_1718; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1720 = 9'hb5 == io_r_req_bits_setIdx ? regs_181_0 : _GEN_1719; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1721 = 9'hb6 == io_r_req_bits_setIdx ? regs_182_0 : _GEN_1720; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1722 = 9'hb7 == io_r_req_bits_setIdx ? regs_183_0 : _GEN_1721; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1723 = 9'hb8 == io_r_req_bits_setIdx ? regs_184_0 : _GEN_1722; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1724 = 9'hb9 == io_r_req_bits_setIdx ? regs_185_0 : _GEN_1723; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1725 = 9'hba == io_r_req_bits_setIdx ? regs_186_0 : _GEN_1724; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1726 = 9'hbb == io_r_req_bits_setIdx ? regs_187_0 : _GEN_1725; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1727 = 9'hbc == io_r_req_bits_setIdx ? regs_188_0 : _GEN_1726; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1728 = 9'hbd == io_r_req_bits_setIdx ? regs_189_0 : _GEN_1727; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1729 = 9'hbe == io_r_req_bits_setIdx ? regs_190_0 : _GEN_1728; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1730 = 9'hbf == io_r_req_bits_setIdx ? regs_191_0 : _GEN_1729; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1731 = 9'hc0 == io_r_req_bits_setIdx ? regs_192_0 : _GEN_1730; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1732 = 9'hc1 == io_r_req_bits_setIdx ? regs_193_0 : _GEN_1731; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1733 = 9'hc2 == io_r_req_bits_setIdx ? regs_194_0 : _GEN_1732; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1734 = 9'hc3 == io_r_req_bits_setIdx ? regs_195_0 : _GEN_1733; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1735 = 9'hc4 == io_r_req_bits_setIdx ? regs_196_0 : _GEN_1734; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1736 = 9'hc5 == io_r_req_bits_setIdx ? regs_197_0 : _GEN_1735; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1737 = 9'hc6 == io_r_req_bits_setIdx ? regs_198_0 : _GEN_1736; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1738 = 9'hc7 == io_r_req_bits_setIdx ? regs_199_0 : _GEN_1737; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1739 = 9'hc8 == io_r_req_bits_setIdx ? regs_200_0 : _GEN_1738; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1740 = 9'hc9 == io_r_req_bits_setIdx ? regs_201_0 : _GEN_1739; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1741 = 9'hca == io_r_req_bits_setIdx ? regs_202_0 : _GEN_1740; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1742 = 9'hcb == io_r_req_bits_setIdx ? regs_203_0 : _GEN_1741; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1743 = 9'hcc == io_r_req_bits_setIdx ? regs_204_0 : _GEN_1742; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1744 = 9'hcd == io_r_req_bits_setIdx ? regs_205_0 : _GEN_1743; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1745 = 9'hce == io_r_req_bits_setIdx ? regs_206_0 : _GEN_1744; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1746 = 9'hcf == io_r_req_bits_setIdx ? regs_207_0 : _GEN_1745; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1747 = 9'hd0 == io_r_req_bits_setIdx ? regs_208_0 : _GEN_1746; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1748 = 9'hd1 == io_r_req_bits_setIdx ? regs_209_0 : _GEN_1747; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1749 = 9'hd2 == io_r_req_bits_setIdx ? regs_210_0 : _GEN_1748; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1750 = 9'hd3 == io_r_req_bits_setIdx ? regs_211_0 : _GEN_1749; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1751 = 9'hd4 == io_r_req_bits_setIdx ? regs_212_0 : _GEN_1750; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1752 = 9'hd5 == io_r_req_bits_setIdx ? regs_213_0 : _GEN_1751; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1753 = 9'hd6 == io_r_req_bits_setIdx ? regs_214_0 : _GEN_1752; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1754 = 9'hd7 == io_r_req_bits_setIdx ? regs_215_0 : _GEN_1753; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1755 = 9'hd8 == io_r_req_bits_setIdx ? regs_216_0 : _GEN_1754; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1756 = 9'hd9 == io_r_req_bits_setIdx ? regs_217_0 : _GEN_1755; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1757 = 9'hda == io_r_req_bits_setIdx ? regs_218_0 : _GEN_1756; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1758 = 9'hdb == io_r_req_bits_setIdx ? regs_219_0 : _GEN_1757; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1759 = 9'hdc == io_r_req_bits_setIdx ? regs_220_0 : _GEN_1758; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1760 = 9'hdd == io_r_req_bits_setIdx ? regs_221_0 : _GEN_1759; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1761 = 9'hde == io_r_req_bits_setIdx ? regs_222_0 : _GEN_1760; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1762 = 9'hdf == io_r_req_bits_setIdx ? regs_223_0 : _GEN_1761; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1763 = 9'he0 == io_r_req_bits_setIdx ? regs_224_0 : _GEN_1762; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1764 = 9'he1 == io_r_req_bits_setIdx ? regs_225_0 : _GEN_1763; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1765 = 9'he2 == io_r_req_bits_setIdx ? regs_226_0 : _GEN_1764; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1766 = 9'he3 == io_r_req_bits_setIdx ? regs_227_0 : _GEN_1765; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1767 = 9'he4 == io_r_req_bits_setIdx ? regs_228_0 : _GEN_1766; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1768 = 9'he5 == io_r_req_bits_setIdx ? regs_229_0 : _GEN_1767; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1769 = 9'he6 == io_r_req_bits_setIdx ? regs_230_0 : _GEN_1768; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1770 = 9'he7 == io_r_req_bits_setIdx ? regs_231_0 : _GEN_1769; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1771 = 9'he8 == io_r_req_bits_setIdx ? regs_232_0 : _GEN_1770; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1772 = 9'he9 == io_r_req_bits_setIdx ? regs_233_0 : _GEN_1771; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1773 = 9'hea == io_r_req_bits_setIdx ? regs_234_0 : _GEN_1772; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1774 = 9'heb == io_r_req_bits_setIdx ? regs_235_0 : _GEN_1773; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1775 = 9'hec == io_r_req_bits_setIdx ? regs_236_0 : _GEN_1774; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1776 = 9'hed == io_r_req_bits_setIdx ? regs_237_0 : _GEN_1775; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1777 = 9'hee == io_r_req_bits_setIdx ? regs_238_0 : _GEN_1776; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1778 = 9'hef == io_r_req_bits_setIdx ? regs_239_0 : _GEN_1777; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1779 = 9'hf0 == io_r_req_bits_setIdx ? regs_240_0 : _GEN_1778; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1780 = 9'hf1 == io_r_req_bits_setIdx ? regs_241_0 : _GEN_1779; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1781 = 9'hf2 == io_r_req_bits_setIdx ? regs_242_0 : _GEN_1780; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1782 = 9'hf3 == io_r_req_bits_setIdx ? regs_243_0 : _GEN_1781; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1783 = 9'hf4 == io_r_req_bits_setIdx ? regs_244_0 : _GEN_1782; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1784 = 9'hf5 == io_r_req_bits_setIdx ? regs_245_0 : _GEN_1783; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1785 = 9'hf6 == io_r_req_bits_setIdx ? regs_246_0 : _GEN_1784; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1786 = 9'hf7 == io_r_req_bits_setIdx ? regs_247_0 : _GEN_1785; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1787 = 9'hf8 == io_r_req_bits_setIdx ? regs_248_0 : _GEN_1786; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1788 = 9'hf9 == io_r_req_bits_setIdx ? regs_249_0 : _GEN_1787; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1789 = 9'hfa == io_r_req_bits_setIdx ? regs_250_0 : _GEN_1788; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1790 = 9'hfb == io_r_req_bits_setIdx ? regs_251_0 : _GEN_1789; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1791 = 9'hfc == io_r_req_bits_setIdx ? regs_252_0 : _GEN_1790; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1792 = 9'hfd == io_r_req_bits_setIdx ? regs_253_0 : _GEN_1791; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1793 = 9'hfe == io_r_req_bits_setIdx ? regs_254_0 : _GEN_1792; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1794 = 9'hff == io_r_req_bits_setIdx ? regs_255_0 : _GEN_1793; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1795 = 9'h100 == io_r_req_bits_setIdx ? regs_256_0 : _GEN_1794; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1796 = 9'h101 == io_r_req_bits_setIdx ? regs_257_0 : _GEN_1795; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1797 = 9'h102 == io_r_req_bits_setIdx ? regs_258_0 : _GEN_1796; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1798 = 9'h103 == io_r_req_bits_setIdx ? regs_259_0 : _GEN_1797; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1799 = 9'h104 == io_r_req_bits_setIdx ? regs_260_0 : _GEN_1798; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1800 = 9'h105 == io_r_req_bits_setIdx ? regs_261_0 : _GEN_1799; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1801 = 9'h106 == io_r_req_bits_setIdx ? regs_262_0 : _GEN_1800; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1802 = 9'h107 == io_r_req_bits_setIdx ? regs_263_0 : _GEN_1801; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1803 = 9'h108 == io_r_req_bits_setIdx ? regs_264_0 : _GEN_1802; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1804 = 9'h109 == io_r_req_bits_setIdx ? regs_265_0 : _GEN_1803; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1805 = 9'h10a == io_r_req_bits_setIdx ? regs_266_0 : _GEN_1804; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1806 = 9'h10b == io_r_req_bits_setIdx ? regs_267_0 : _GEN_1805; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1807 = 9'h10c == io_r_req_bits_setIdx ? regs_268_0 : _GEN_1806; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1808 = 9'h10d == io_r_req_bits_setIdx ? regs_269_0 : _GEN_1807; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1809 = 9'h10e == io_r_req_bits_setIdx ? regs_270_0 : _GEN_1808; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1810 = 9'h10f == io_r_req_bits_setIdx ? regs_271_0 : _GEN_1809; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1811 = 9'h110 == io_r_req_bits_setIdx ? regs_272_0 : _GEN_1810; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1812 = 9'h111 == io_r_req_bits_setIdx ? regs_273_0 : _GEN_1811; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1813 = 9'h112 == io_r_req_bits_setIdx ? regs_274_0 : _GEN_1812; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1814 = 9'h113 == io_r_req_bits_setIdx ? regs_275_0 : _GEN_1813; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1815 = 9'h114 == io_r_req_bits_setIdx ? regs_276_0 : _GEN_1814; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1816 = 9'h115 == io_r_req_bits_setIdx ? regs_277_0 : _GEN_1815; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1817 = 9'h116 == io_r_req_bits_setIdx ? regs_278_0 : _GEN_1816; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1818 = 9'h117 == io_r_req_bits_setIdx ? regs_279_0 : _GEN_1817; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1819 = 9'h118 == io_r_req_bits_setIdx ? regs_280_0 : _GEN_1818; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1820 = 9'h119 == io_r_req_bits_setIdx ? regs_281_0 : _GEN_1819; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1821 = 9'h11a == io_r_req_bits_setIdx ? regs_282_0 : _GEN_1820; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1822 = 9'h11b == io_r_req_bits_setIdx ? regs_283_0 : _GEN_1821; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1823 = 9'h11c == io_r_req_bits_setIdx ? regs_284_0 : _GEN_1822; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1824 = 9'h11d == io_r_req_bits_setIdx ? regs_285_0 : _GEN_1823; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1825 = 9'h11e == io_r_req_bits_setIdx ? regs_286_0 : _GEN_1824; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1826 = 9'h11f == io_r_req_bits_setIdx ? regs_287_0 : _GEN_1825; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1827 = 9'h120 == io_r_req_bits_setIdx ? regs_288_0 : _GEN_1826; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1828 = 9'h121 == io_r_req_bits_setIdx ? regs_289_0 : _GEN_1827; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1829 = 9'h122 == io_r_req_bits_setIdx ? regs_290_0 : _GEN_1828; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1830 = 9'h123 == io_r_req_bits_setIdx ? regs_291_0 : _GEN_1829; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1831 = 9'h124 == io_r_req_bits_setIdx ? regs_292_0 : _GEN_1830; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1832 = 9'h125 == io_r_req_bits_setIdx ? regs_293_0 : _GEN_1831; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1833 = 9'h126 == io_r_req_bits_setIdx ? regs_294_0 : _GEN_1832; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1834 = 9'h127 == io_r_req_bits_setIdx ? regs_295_0 : _GEN_1833; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1835 = 9'h128 == io_r_req_bits_setIdx ? regs_296_0 : _GEN_1834; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1836 = 9'h129 == io_r_req_bits_setIdx ? regs_297_0 : _GEN_1835; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1837 = 9'h12a == io_r_req_bits_setIdx ? regs_298_0 : _GEN_1836; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1838 = 9'h12b == io_r_req_bits_setIdx ? regs_299_0 : _GEN_1837; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1839 = 9'h12c == io_r_req_bits_setIdx ? regs_300_0 : _GEN_1838; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1840 = 9'h12d == io_r_req_bits_setIdx ? regs_301_0 : _GEN_1839; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1841 = 9'h12e == io_r_req_bits_setIdx ? regs_302_0 : _GEN_1840; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1842 = 9'h12f == io_r_req_bits_setIdx ? regs_303_0 : _GEN_1841; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1843 = 9'h130 == io_r_req_bits_setIdx ? regs_304_0 : _GEN_1842; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1844 = 9'h131 == io_r_req_bits_setIdx ? regs_305_0 : _GEN_1843; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1845 = 9'h132 == io_r_req_bits_setIdx ? regs_306_0 : _GEN_1844; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1846 = 9'h133 == io_r_req_bits_setIdx ? regs_307_0 : _GEN_1845; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1847 = 9'h134 == io_r_req_bits_setIdx ? regs_308_0 : _GEN_1846; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1848 = 9'h135 == io_r_req_bits_setIdx ? regs_309_0 : _GEN_1847; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1849 = 9'h136 == io_r_req_bits_setIdx ? regs_310_0 : _GEN_1848; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1850 = 9'h137 == io_r_req_bits_setIdx ? regs_311_0 : _GEN_1849; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1851 = 9'h138 == io_r_req_bits_setIdx ? regs_312_0 : _GEN_1850; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1852 = 9'h139 == io_r_req_bits_setIdx ? regs_313_0 : _GEN_1851; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1853 = 9'h13a == io_r_req_bits_setIdx ? regs_314_0 : _GEN_1852; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1854 = 9'h13b == io_r_req_bits_setIdx ? regs_315_0 : _GEN_1853; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1855 = 9'h13c == io_r_req_bits_setIdx ? regs_316_0 : _GEN_1854; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1856 = 9'h13d == io_r_req_bits_setIdx ? regs_317_0 : _GEN_1855; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1857 = 9'h13e == io_r_req_bits_setIdx ? regs_318_0 : _GEN_1856; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1858 = 9'h13f == io_r_req_bits_setIdx ? regs_319_0 : _GEN_1857; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1859 = 9'h140 == io_r_req_bits_setIdx ? regs_320_0 : _GEN_1858; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1860 = 9'h141 == io_r_req_bits_setIdx ? regs_321_0 : _GEN_1859; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1861 = 9'h142 == io_r_req_bits_setIdx ? regs_322_0 : _GEN_1860; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1862 = 9'h143 == io_r_req_bits_setIdx ? regs_323_0 : _GEN_1861; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1863 = 9'h144 == io_r_req_bits_setIdx ? regs_324_0 : _GEN_1862; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1864 = 9'h145 == io_r_req_bits_setIdx ? regs_325_0 : _GEN_1863; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1865 = 9'h146 == io_r_req_bits_setIdx ? regs_326_0 : _GEN_1864; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1866 = 9'h147 == io_r_req_bits_setIdx ? regs_327_0 : _GEN_1865; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1867 = 9'h148 == io_r_req_bits_setIdx ? regs_328_0 : _GEN_1866; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1868 = 9'h149 == io_r_req_bits_setIdx ? regs_329_0 : _GEN_1867; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1869 = 9'h14a == io_r_req_bits_setIdx ? regs_330_0 : _GEN_1868; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1870 = 9'h14b == io_r_req_bits_setIdx ? regs_331_0 : _GEN_1869; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1871 = 9'h14c == io_r_req_bits_setIdx ? regs_332_0 : _GEN_1870; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1872 = 9'h14d == io_r_req_bits_setIdx ? regs_333_0 : _GEN_1871; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1873 = 9'h14e == io_r_req_bits_setIdx ? regs_334_0 : _GEN_1872; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1874 = 9'h14f == io_r_req_bits_setIdx ? regs_335_0 : _GEN_1873; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1875 = 9'h150 == io_r_req_bits_setIdx ? regs_336_0 : _GEN_1874; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1876 = 9'h151 == io_r_req_bits_setIdx ? regs_337_0 : _GEN_1875; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1877 = 9'h152 == io_r_req_bits_setIdx ? regs_338_0 : _GEN_1876; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1878 = 9'h153 == io_r_req_bits_setIdx ? regs_339_0 : _GEN_1877; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1879 = 9'h154 == io_r_req_bits_setIdx ? regs_340_0 : _GEN_1878; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1880 = 9'h155 == io_r_req_bits_setIdx ? regs_341_0 : _GEN_1879; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1881 = 9'h156 == io_r_req_bits_setIdx ? regs_342_0 : _GEN_1880; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1882 = 9'h157 == io_r_req_bits_setIdx ? regs_343_0 : _GEN_1881; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1883 = 9'h158 == io_r_req_bits_setIdx ? regs_344_0 : _GEN_1882; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1884 = 9'h159 == io_r_req_bits_setIdx ? regs_345_0 : _GEN_1883; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1885 = 9'h15a == io_r_req_bits_setIdx ? regs_346_0 : _GEN_1884; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1886 = 9'h15b == io_r_req_bits_setIdx ? regs_347_0 : _GEN_1885; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1887 = 9'h15c == io_r_req_bits_setIdx ? regs_348_0 : _GEN_1886; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1888 = 9'h15d == io_r_req_bits_setIdx ? regs_349_0 : _GEN_1887; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1889 = 9'h15e == io_r_req_bits_setIdx ? regs_350_0 : _GEN_1888; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1890 = 9'h15f == io_r_req_bits_setIdx ? regs_351_0 : _GEN_1889; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1891 = 9'h160 == io_r_req_bits_setIdx ? regs_352_0 : _GEN_1890; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1892 = 9'h161 == io_r_req_bits_setIdx ? regs_353_0 : _GEN_1891; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1893 = 9'h162 == io_r_req_bits_setIdx ? regs_354_0 : _GEN_1892; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1894 = 9'h163 == io_r_req_bits_setIdx ? regs_355_0 : _GEN_1893; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1895 = 9'h164 == io_r_req_bits_setIdx ? regs_356_0 : _GEN_1894; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1896 = 9'h165 == io_r_req_bits_setIdx ? regs_357_0 : _GEN_1895; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1897 = 9'h166 == io_r_req_bits_setIdx ? regs_358_0 : _GEN_1896; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1898 = 9'h167 == io_r_req_bits_setIdx ? regs_359_0 : _GEN_1897; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1899 = 9'h168 == io_r_req_bits_setIdx ? regs_360_0 : _GEN_1898; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1900 = 9'h169 == io_r_req_bits_setIdx ? regs_361_0 : _GEN_1899; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1901 = 9'h16a == io_r_req_bits_setIdx ? regs_362_0 : _GEN_1900; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1902 = 9'h16b == io_r_req_bits_setIdx ? regs_363_0 : _GEN_1901; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1903 = 9'h16c == io_r_req_bits_setIdx ? regs_364_0 : _GEN_1902; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1904 = 9'h16d == io_r_req_bits_setIdx ? regs_365_0 : _GEN_1903; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1905 = 9'h16e == io_r_req_bits_setIdx ? regs_366_0 : _GEN_1904; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1906 = 9'h16f == io_r_req_bits_setIdx ? regs_367_0 : _GEN_1905; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1907 = 9'h170 == io_r_req_bits_setIdx ? regs_368_0 : _GEN_1906; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1908 = 9'h171 == io_r_req_bits_setIdx ? regs_369_0 : _GEN_1907; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1909 = 9'h172 == io_r_req_bits_setIdx ? regs_370_0 : _GEN_1908; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1910 = 9'h173 == io_r_req_bits_setIdx ? regs_371_0 : _GEN_1909; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1911 = 9'h174 == io_r_req_bits_setIdx ? regs_372_0 : _GEN_1910; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1912 = 9'h175 == io_r_req_bits_setIdx ? regs_373_0 : _GEN_1911; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1913 = 9'h176 == io_r_req_bits_setIdx ? regs_374_0 : _GEN_1912; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1914 = 9'h177 == io_r_req_bits_setIdx ? regs_375_0 : _GEN_1913; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1915 = 9'h178 == io_r_req_bits_setIdx ? regs_376_0 : _GEN_1914; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1916 = 9'h179 == io_r_req_bits_setIdx ? regs_377_0 : _GEN_1915; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1917 = 9'h17a == io_r_req_bits_setIdx ? regs_378_0 : _GEN_1916; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1918 = 9'h17b == io_r_req_bits_setIdx ? regs_379_0 : _GEN_1917; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1919 = 9'h17c == io_r_req_bits_setIdx ? regs_380_0 : _GEN_1918; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1920 = 9'h17d == io_r_req_bits_setIdx ? regs_381_0 : _GEN_1919; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1921 = 9'h17e == io_r_req_bits_setIdx ? regs_382_0 : _GEN_1920; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1922 = 9'h17f == io_r_req_bits_setIdx ? regs_383_0 : _GEN_1921; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1923 = 9'h180 == io_r_req_bits_setIdx ? regs_384_0 : _GEN_1922; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1924 = 9'h181 == io_r_req_bits_setIdx ? regs_385_0 : _GEN_1923; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1925 = 9'h182 == io_r_req_bits_setIdx ? regs_386_0 : _GEN_1924; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1926 = 9'h183 == io_r_req_bits_setIdx ? regs_387_0 : _GEN_1925; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1927 = 9'h184 == io_r_req_bits_setIdx ? regs_388_0 : _GEN_1926; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1928 = 9'h185 == io_r_req_bits_setIdx ? regs_389_0 : _GEN_1927; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1929 = 9'h186 == io_r_req_bits_setIdx ? regs_390_0 : _GEN_1928; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1930 = 9'h187 == io_r_req_bits_setIdx ? regs_391_0 : _GEN_1929; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1931 = 9'h188 == io_r_req_bits_setIdx ? regs_392_0 : _GEN_1930; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1932 = 9'h189 == io_r_req_bits_setIdx ? regs_393_0 : _GEN_1931; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1933 = 9'h18a == io_r_req_bits_setIdx ? regs_394_0 : _GEN_1932; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1934 = 9'h18b == io_r_req_bits_setIdx ? regs_395_0 : _GEN_1933; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1935 = 9'h18c == io_r_req_bits_setIdx ? regs_396_0 : _GEN_1934; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1936 = 9'h18d == io_r_req_bits_setIdx ? regs_397_0 : _GEN_1935; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1937 = 9'h18e == io_r_req_bits_setIdx ? regs_398_0 : _GEN_1936; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1938 = 9'h18f == io_r_req_bits_setIdx ? regs_399_0 : _GEN_1937; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1939 = 9'h190 == io_r_req_bits_setIdx ? regs_400_0 : _GEN_1938; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1940 = 9'h191 == io_r_req_bits_setIdx ? regs_401_0 : _GEN_1939; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1941 = 9'h192 == io_r_req_bits_setIdx ? regs_402_0 : _GEN_1940; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1942 = 9'h193 == io_r_req_bits_setIdx ? regs_403_0 : _GEN_1941; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1943 = 9'h194 == io_r_req_bits_setIdx ? regs_404_0 : _GEN_1942; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1944 = 9'h195 == io_r_req_bits_setIdx ? regs_405_0 : _GEN_1943; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1945 = 9'h196 == io_r_req_bits_setIdx ? regs_406_0 : _GEN_1944; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1946 = 9'h197 == io_r_req_bits_setIdx ? regs_407_0 : _GEN_1945; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1947 = 9'h198 == io_r_req_bits_setIdx ? regs_408_0 : _GEN_1946; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1948 = 9'h199 == io_r_req_bits_setIdx ? regs_409_0 : _GEN_1947; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1949 = 9'h19a == io_r_req_bits_setIdx ? regs_410_0 : _GEN_1948; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1950 = 9'h19b == io_r_req_bits_setIdx ? regs_411_0 : _GEN_1949; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1951 = 9'h19c == io_r_req_bits_setIdx ? regs_412_0 : _GEN_1950; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1952 = 9'h19d == io_r_req_bits_setIdx ? regs_413_0 : _GEN_1951; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1953 = 9'h19e == io_r_req_bits_setIdx ? regs_414_0 : _GEN_1952; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1954 = 9'h19f == io_r_req_bits_setIdx ? regs_415_0 : _GEN_1953; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1955 = 9'h1a0 == io_r_req_bits_setIdx ? regs_416_0 : _GEN_1954; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1956 = 9'h1a1 == io_r_req_bits_setIdx ? regs_417_0 : _GEN_1955; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1957 = 9'h1a2 == io_r_req_bits_setIdx ? regs_418_0 : _GEN_1956; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1958 = 9'h1a3 == io_r_req_bits_setIdx ? regs_419_0 : _GEN_1957; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1959 = 9'h1a4 == io_r_req_bits_setIdx ? regs_420_0 : _GEN_1958; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1960 = 9'h1a5 == io_r_req_bits_setIdx ? regs_421_0 : _GEN_1959; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1961 = 9'h1a6 == io_r_req_bits_setIdx ? regs_422_0 : _GEN_1960; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1962 = 9'h1a7 == io_r_req_bits_setIdx ? regs_423_0 : _GEN_1961; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1963 = 9'h1a8 == io_r_req_bits_setIdx ? regs_424_0 : _GEN_1962; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1964 = 9'h1a9 == io_r_req_bits_setIdx ? regs_425_0 : _GEN_1963; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1965 = 9'h1aa == io_r_req_bits_setIdx ? regs_426_0 : _GEN_1964; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1966 = 9'h1ab == io_r_req_bits_setIdx ? regs_427_0 : _GEN_1965; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1967 = 9'h1ac == io_r_req_bits_setIdx ? regs_428_0 : _GEN_1966; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1968 = 9'h1ad == io_r_req_bits_setIdx ? regs_429_0 : _GEN_1967; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1969 = 9'h1ae == io_r_req_bits_setIdx ? regs_430_0 : _GEN_1968; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1970 = 9'h1af == io_r_req_bits_setIdx ? regs_431_0 : _GEN_1969; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1971 = 9'h1b0 == io_r_req_bits_setIdx ? regs_432_0 : _GEN_1970; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1972 = 9'h1b1 == io_r_req_bits_setIdx ? regs_433_0 : _GEN_1971; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1973 = 9'h1b2 == io_r_req_bits_setIdx ? regs_434_0 : _GEN_1972; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1974 = 9'h1b3 == io_r_req_bits_setIdx ? regs_435_0 : _GEN_1973; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1975 = 9'h1b4 == io_r_req_bits_setIdx ? regs_436_0 : _GEN_1974; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1976 = 9'h1b5 == io_r_req_bits_setIdx ? regs_437_0 : _GEN_1975; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1977 = 9'h1b6 == io_r_req_bits_setIdx ? regs_438_0 : _GEN_1976; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1978 = 9'h1b7 == io_r_req_bits_setIdx ? regs_439_0 : _GEN_1977; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1979 = 9'h1b8 == io_r_req_bits_setIdx ? regs_440_0 : _GEN_1978; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1980 = 9'h1b9 == io_r_req_bits_setIdx ? regs_441_0 : _GEN_1979; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1981 = 9'h1ba == io_r_req_bits_setIdx ? regs_442_0 : _GEN_1980; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1982 = 9'h1bb == io_r_req_bits_setIdx ? regs_443_0 : _GEN_1981; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1983 = 9'h1bc == io_r_req_bits_setIdx ? regs_444_0 : _GEN_1982; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1984 = 9'h1bd == io_r_req_bits_setIdx ? regs_445_0 : _GEN_1983; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1985 = 9'h1be == io_r_req_bits_setIdx ? regs_446_0 : _GEN_1984; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1986 = 9'h1bf == io_r_req_bits_setIdx ? regs_447_0 : _GEN_1985; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1987 = 9'h1c0 == io_r_req_bits_setIdx ? regs_448_0 : _GEN_1986; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1988 = 9'h1c1 == io_r_req_bits_setIdx ? regs_449_0 : _GEN_1987; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1989 = 9'h1c2 == io_r_req_bits_setIdx ? regs_450_0 : _GEN_1988; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1990 = 9'h1c3 == io_r_req_bits_setIdx ? regs_451_0 : _GEN_1989; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1991 = 9'h1c4 == io_r_req_bits_setIdx ? regs_452_0 : _GEN_1990; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1992 = 9'h1c5 == io_r_req_bits_setIdx ? regs_453_0 : _GEN_1991; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1993 = 9'h1c6 == io_r_req_bits_setIdx ? regs_454_0 : _GEN_1992; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1994 = 9'h1c7 == io_r_req_bits_setIdx ? regs_455_0 : _GEN_1993; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1995 = 9'h1c8 == io_r_req_bits_setIdx ? regs_456_0 : _GEN_1994; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1996 = 9'h1c9 == io_r_req_bits_setIdx ? regs_457_0 : _GEN_1995; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1997 = 9'h1ca == io_r_req_bits_setIdx ? regs_458_0 : _GEN_1996; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1998 = 9'h1cb == io_r_req_bits_setIdx ? regs_459_0 : _GEN_1997; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_1999 = 9'h1cc == io_r_req_bits_setIdx ? regs_460_0 : _GEN_1998; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2000 = 9'h1cd == io_r_req_bits_setIdx ? regs_461_0 : _GEN_1999; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2001 = 9'h1ce == io_r_req_bits_setIdx ? regs_462_0 : _GEN_2000; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2002 = 9'h1cf == io_r_req_bits_setIdx ? regs_463_0 : _GEN_2001; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2003 = 9'h1d0 == io_r_req_bits_setIdx ? regs_464_0 : _GEN_2002; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2004 = 9'h1d1 == io_r_req_bits_setIdx ? regs_465_0 : _GEN_2003; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2005 = 9'h1d2 == io_r_req_bits_setIdx ? regs_466_0 : _GEN_2004; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2006 = 9'h1d3 == io_r_req_bits_setIdx ? regs_467_0 : _GEN_2005; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2007 = 9'h1d4 == io_r_req_bits_setIdx ? regs_468_0 : _GEN_2006; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2008 = 9'h1d5 == io_r_req_bits_setIdx ? regs_469_0 : _GEN_2007; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2009 = 9'h1d6 == io_r_req_bits_setIdx ? regs_470_0 : _GEN_2008; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2010 = 9'h1d7 == io_r_req_bits_setIdx ? regs_471_0 : _GEN_2009; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2011 = 9'h1d8 == io_r_req_bits_setIdx ? regs_472_0 : _GEN_2010; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2012 = 9'h1d9 == io_r_req_bits_setIdx ? regs_473_0 : _GEN_2011; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2013 = 9'h1da == io_r_req_bits_setIdx ? regs_474_0 : _GEN_2012; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2014 = 9'h1db == io_r_req_bits_setIdx ? regs_475_0 : _GEN_2013; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2015 = 9'h1dc == io_r_req_bits_setIdx ? regs_476_0 : _GEN_2014; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2016 = 9'h1dd == io_r_req_bits_setIdx ? regs_477_0 : _GEN_2015; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2017 = 9'h1de == io_r_req_bits_setIdx ? regs_478_0 : _GEN_2016; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2018 = 9'h1df == io_r_req_bits_setIdx ? regs_479_0 : _GEN_2017; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2019 = 9'h1e0 == io_r_req_bits_setIdx ? regs_480_0 : _GEN_2018; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2020 = 9'h1e1 == io_r_req_bits_setIdx ? regs_481_0 : _GEN_2019; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2021 = 9'h1e2 == io_r_req_bits_setIdx ? regs_482_0 : _GEN_2020; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2022 = 9'h1e3 == io_r_req_bits_setIdx ? regs_483_0 : _GEN_2021; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2023 = 9'h1e4 == io_r_req_bits_setIdx ? regs_484_0 : _GEN_2022; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2024 = 9'h1e5 == io_r_req_bits_setIdx ? regs_485_0 : _GEN_2023; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2025 = 9'h1e6 == io_r_req_bits_setIdx ? regs_486_0 : _GEN_2024; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2026 = 9'h1e7 == io_r_req_bits_setIdx ? regs_487_0 : _GEN_2025; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2027 = 9'h1e8 == io_r_req_bits_setIdx ? regs_488_0 : _GEN_2026; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2028 = 9'h1e9 == io_r_req_bits_setIdx ? regs_489_0 : _GEN_2027; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2029 = 9'h1ea == io_r_req_bits_setIdx ? regs_490_0 : _GEN_2028; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2030 = 9'h1eb == io_r_req_bits_setIdx ? regs_491_0 : _GEN_2029; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2031 = 9'h1ec == io_r_req_bits_setIdx ? regs_492_0 : _GEN_2030; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2032 = 9'h1ed == io_r_req_bits_setIdx ? regs_493_0 : _GEN_2031; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2033 = 9'h1ee == io_r_req_bits_setIdx ? regs_494_0 : _GEN_2032; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2034 = 9'h1ef == io_r_req_bits_setIdx ? regs_495_0 : _GEN_2033; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2035 = 9'h1f0 == io_r_req_bits_setIdx ? regs_496_0 : _GEN_2034; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2036 = 9'h1f1 == io_r_req_bits_setIdx ? regs_497_0 : _GEN_2035; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2037 = 9'h1f2 == io_r_req_bits_setIdx ? regs_498_0 : _GEN_2036; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2038 = 9'h1f3 == io_r_req_bits_setIdx ? regs_499_0 : _GEN_2037; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2039 = 9'h1f4 == io_r_req_bits_setIdx ? regs_500_0 : _GEN_2038; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2040 = 9'h1f5 == io_r_req_bits_setIdx ? regs_501_0 : _GEN_2039; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2041 = 9'h1f6 == io_r_req_bits_setIdx ? regs_502_0 : _GEN_2040; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2042 = 9'h1f7 == io_r_req_bits_setIdx ? regs_503_0 : _GEN_2041; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2043 = 9'h1f8 == io_r_req_bits_setIdx ? regs_504_0 : _GEN_2042; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2044 = 9'h1f9 == io_r_req_bits_setIdx ? regs_505_0 : _GEN_2043; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2045 = 9'h1fa == io_r_req_bits_setIdx ? regs_506_0 : _GEN_2044; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2046 = 9'h1fb == io_r_req_bits_setIdx ? regs_507_0 : _GEN_2045; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  wire [72:0] _GEN_2047 = 9'h1fc == io_r_req_bits_setIdx ? regs_508_0 : _GEN_2046; // @[src/main/scala/utils/RegMem.scala 39:{14,14}]
  reg  rdata_REG; // @[src/main/scala/utils/Hold.scala 29:110]
  reg [72:0] rdata_r_1_0; // @[src/main/scala/utils/Hold.scala 23:65]
  wire [72:0] _GEN_2052 = rdata_REG ? rdata_r_0 : rdata_r_1_0; // @[src/main/scala/utils/Hold.scala 23:{65,65,65}]
  assign io_r_req_ready = ~resetState & _realRen_T; // @[src/main/scala/utils/SRAMTemplate.scala 101:33]
  assign io_r_resp_data_0_tag = _GEN_2052[72:45]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign io_r_resp_data_0__type = _GEN_2052[44:43]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign io_r_resp_data_0_target = _GEN_2052[42:4]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign io_r_resp_data_0_brIdx = _GEN_2052[3:1]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign io_r_resp_data_0_valid = _GEN_2052[0]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_0_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h0 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_0_0 <= 73'h0;
        end else begin
          regs_0_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_1_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_1_0 <= 73'h0;
        end else begin
          regs_1_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_2_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h2 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_2_0 <= 73'h0;
        end else begin
          regs_2_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_3_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h3 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_3_0 <= 73'h0;
        end else begin
          regs_3_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_4_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h4 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_4_0 <= 73'h0;
        end else begin
          regs_4_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_5_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h5 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_5_0 <= 73'h0;
        end else begin
          regs_5_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_6_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h6 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_6_0 <= 73'h0;
        end else begin
          regs_6_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_7_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h7 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_7_0 <= 73'h0;
        end else begin
          regs_7_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_8_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h8 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_8_0 <= 73'h0;
        end else begin
          regs_8_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_9_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h9 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_9_0 <= 73'h0;
        end else begin
          regs_9_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_10_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'ha == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_10_0 <= 73'h0;
        end else begin
          regs_10_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_11_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hb == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_11_0 <= 73'h0;
        end else begin
          regs_11_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_12_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hc == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_12_0 <= 73'h0;
        end else begin
          regs_12_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_13_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hd == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_13_0 <= 73'h0;
        end else begin
          regs_13_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_14_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'he == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_14_0 <= 73'h0;
        end else begin
          regs_14_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_15_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hf == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_15_0 <= 73'h0;
        end else begin
          regs_15_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_16_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h10 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_16_0 <= 73'h0;
        end else begin
          regs_16_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_17_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h11 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_17_0 <= 73'h0;
        end else begin
          regs_17_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_18_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h12 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_18_0 <= 73'h0;
        end else begin
          regs_18_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_19_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h13 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_19_0 <= 73'h0;
        end else begin
          regs_19_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_20_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h14 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_20_0 <= 73'h0;
        end else begin
          regs_20_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_21_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h15 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_21_0 <= 73'h0;
        end else begin
          regs_21_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_22_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h16 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_22_0 <= 73'h0;
        end else begin
          regs_22_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_23_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h17 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_23_0 <= 73'h0;
        end else begin
          regs_23_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_24_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h18 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_24_0 <= 73'h0;
        end else begin
          regs_24_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_25_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h19 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_25_0 <= 73'h0;
        end else begin
          regs_25_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_26_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1a == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_26_0 <= 73'h0;
        end else begin
          regs_26_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_27_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1b == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_27_0 <= 73'h0;
        end else begin
          regs_27_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_28_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1c == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_28_0 <= 73'h0;
        end else begin
          regs_28_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_29_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1d == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_29_0 <= 73'h0;
        end else begin
          regs_29_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_30_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1e == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_30_0 <= 73'h0;
        end else begin
          regs_30_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_31_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1f == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_31_0 <= 73'h0;
        end else begin
          regs_31_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_32_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h20 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_32_0 <= 73'h0;
        end else begin
          regs_32_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_33_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h21 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_33_0 <= 73'h0;
        end else begin
          regs_33_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_34_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h22 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_34_0 <= 73'h0;
        end else begin
          regs_34_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_35_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h23 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_35_0 <= 73'h0;
        end else begin
          regs_35_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_36_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h24 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_36_0 <= 73'h0;
        end else begin
          regs_36_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_37_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h25 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_37_0 <= 73'h0;
        end else begin
          regs_37_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_38_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h26 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_38_0 <= 73'h0;
        end else begin
          regs_38_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_39_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h27 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_39_0 <= 73'h0;
        end else begin
          regs_39_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_40_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h28 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_40_0 <= 73'h0;
        end else begin
          regs_40_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_41_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h29 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_41_0 <= 73'h0;
        end else begin
          regs_41_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_42_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h2a == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_42_0 <= 73'h0;
        end else begin
          regs_42_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_43_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h2b == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_43_0 <= 73'h0;
        end else begin
          regs_43_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_44_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h2c == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_44_0 <= 73'h0;
        end else begin
          regs_44_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_45_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h2d == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_45_0 <= 73'h0;
        end else begin
          regs_45_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_46_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h2e == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_46_0 <= 73'h0;
        end else begin
          regs_46_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_47_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h2f == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_47_0 <= 73'h0;
        end else begin
          regs_47_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_48_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h30 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_48_0 <= 73'h0;
        end else begin
          regs_48_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_49_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h31 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_49_0 <= 73'h0;
        end else begin
          regs_49_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_50_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h32 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_50_0 <= 73'h0;
        end else begin
          regs_50_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_51_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h33 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_51_0 <= 73'h0;
        end else begin
          regs_51_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_52_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h34 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_52_0 <= 73'h0;
        end else begin
          regs_52_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_53_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h35 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_53_0 <= 73'h0;
        end else begin
          regs_53_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_54_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h36 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_54_0 <= 73'h0;
        end else begin
          regs_54_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_55_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h37 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_55_0 <= 73'h0;
        end else begin
          regs_55_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_56_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h38 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_56_0 <= 73'h0;
        end else begin
          regs_56_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_57_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h39 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_57_0 <= 73'h0;
        end else begin
          regs_57_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_58_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h3a == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_58_0 <= 73'h0;
        end else begin
          regs_58_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_59_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h3b == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_59_0 <= 73'h0;
        end else begin
          regs_59_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_60_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h3c == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_60_0 <= 73'h0;
        end else begin
          regs_60_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_61_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h3d == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_61_0 <= 73'h0;
        end else begin
          regs_61_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_62_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h3e == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_62_0 <= 73'h0;
        end else begin
          regs_62_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_63_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h3f == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_63_0 <= 73'h0;
        end else begin
          regs_63_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_64_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h40 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_64_0 <= 73'h0;
        end else begin
          regs_64_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_65_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h41 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_65_0 <= 73'h0;
        end else begin
          regs_65_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_66_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h42 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_66_0 <= 73'h0;
        end else begin
          regs_66_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_67_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h43 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_67_0 <= 73'h0;
        end else begin
          regs_67_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_68_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h44 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_68_0 <= 73'h0;
        end else begin
          regs_68_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_69_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h45 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_69_0 <= 73'h0;
        end else begin
          regs_69_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_70_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h46 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_70_0 <= 73'h0;
        end else begin
          regs_70_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_71_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h47 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_71_0 <= 73'h0;
        end else begin
          regs_71_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_72_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h48 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_72_0 <= 73'h0;
        end else begin
          regs_72_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_73_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h49 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_73_0 <= 73'h0;
        end else begin
          regs_73_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_74_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h4a == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_74_0 <= 73'h0;
        end else begin
          regs_74_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_75_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h4b == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_75_0 <= 73'h0;
        end else begin
          regs_75_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_76_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h4c == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_76_0 <= 73'h0;
        end else begin
          regs_76_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_77_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h4d == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_77_0 <= 73'h0;
        end else begin
          regs_77_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_78_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h4e == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_78_0 <= 73'h0;
        end else begin
          regs_78_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_79_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h4f == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_79_0 <= 73'h0;
        end else begin
          regs_79_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_80_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h50 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_80_0 <= 73'h0;
        end else begin
          regs_80_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_81_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h51 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_81_0 <= 73'h0;
        end else begin
          regs_81_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_82_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h52 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_82_0 <= 73'h0;
        end else begin
          regs_82_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_83_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h53 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_83_0 <= 73'h0;
        end else begin
          regs_83_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_84_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h54 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_84_0 <= 73'h0;
        end else begin
          regs_84_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_85_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h55 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_85_0 <= 73'h0;
        end else begin
          regs_85_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_86_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h56 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_86_0 <= 73'h0;
        end else begin
          regs_86_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_87_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h57 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_87_0 <= 73'h0;
        end else begin
          regs_87_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_88_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h58 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_88_0 <= 73'h0;
        end else begin
          regs_88_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_89_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h59 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_89_0 <= 73'h0;
        end else begin
          regs_89_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_90_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h5a == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_90_0 <= 73'h0;
        end else begin
          regs_90_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_91_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h5b == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_91_0 <= 73'h0;
        end else begin
          regs_91_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_92_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h5c == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_92_0 <= 73'h0;
        end else begin
          regs_92_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_93_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h5d == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_93_0 <= 73'h0;
        end else begin
          regs_93_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_94_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h5e == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_94_0 <= 73'h0;
        end else begin
          regs_94_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_95_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h5f == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_95_0 <= 73'h0;
        end else begin
          regs_95_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_96_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h60 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_96_0 <= 73'h0;
        end else begin
          regs_96_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_97_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h61 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_97_0 <= 73'h0;
        end else begin
          regs_97_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_98_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h62 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_98_0 <= 73'h0;
        end else begin
          regs_98_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_99_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h63 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_99_0 <= 73'h0;
        end else begin
          regs_99_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_100_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h64 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_100_0 <= 73'h0;
        end else begin
          regs_100_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_101_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h65 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_101_0 <= 73'h0;
        end else begin
          regs_101_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_102_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h66 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_102_0 <= 73'h0;
        end else begin
          regs_102_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_103_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h67 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_103_0 <= 73'h0;
        end else begin
          regs_103_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_104_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h68 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_104_0 <= 73'h0;
        end else begin
          regs_104_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_105_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h69 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_105_0 <= 73'h0;
        end else begin
          regs_105_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_106_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h6a == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_106_0 <= 73'h0;
        end else begin
          regs_106_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_107_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h6b == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_107_0 <= 73'h0;
        end else begin
          regs_107_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_108_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h6c == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_108_0 <= 73'h0;
        end else begin
          regs_108_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_109_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h6d == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_109_0 <= 73'h0;
        end else begin
          regs_109_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_110_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h6e == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_110_0 <= 73'h0;
        end else begin
          regs_110_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_111_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h6f == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_111_0 <= 73'h0;
        end else begin
          regs_111_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_112_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h70 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_112_0 <= 73'h0;
        end else begin
          regs_112_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_113_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h71 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_113_0 <= 73'h0;
        end else begin
          regs_113_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_114_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h72 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_114_0 <= 73'h0;
        end else begin
          regs_114_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_115_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h73 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_115_0 <= 73'h0;
        end else begin
          regs_115_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_116_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h74 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_116_0 <= 73'h0;
        end else begin
          regs_116_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_117_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h75 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_117_0 <= 73'h0;
        end else begin
          regs_117_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_118_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h76 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_118_0 <= 73'h0;
        end else begin
          regs_118_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_119_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h77 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_119_0 <= 73'h0;
        end else begin
          regs_119_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_120_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h78 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_120_0 <= 73'h0;
        end else begin
          regs_120_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_121_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h79 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_121_0 <= 73'h0;
        end else begin
          regs_121_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_122_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h7a == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_122_0 <= 73'h0;
        end else begin
          regs_122_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_123_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h7b == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_123_0 <= 73'h0;
        end else begin
          regs_123_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_124_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h7c == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_124_0 <= 73'h0;
        end else begin
          regs_124_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_125_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h7d == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_125_0 <= 73'h0;
        end else begin
          regs_125_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_126_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h7e == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_126_0 <= 73'h0;
        end else begin
          regs_126_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_127_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h7f == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_127_0 <= 73'h0;
        end else begin
          regs_127_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_128_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h80 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_128_0 <= 73'h0;
        end else begin
          regs_128_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_129_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h81 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_129_0 <= 73'h0;
        end else begin
          regs_129_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_130_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h82 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_130_0 <= 73'h0;
        end else begin
          regs_130_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_131_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h83 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_131_0 <= 73'h0;
        end else begin
          regs_131_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_132_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h84 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_132_0 <= 73'h0;
        end else begin
          regs_132_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_133_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h85 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_133_0 <= 73'h0;
        end else begin
          regs_133_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_134_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h86 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_134_0 <= 73'h0;
        end else begin
          regs_134_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_135_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h87 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_135_0 <= 73'h0;
        end else begin
          regs_135_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_136_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h88 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_136_0 <= 73'h0;
        end else begin
          regs_136_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_137_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h89 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_137_0 <= 73'h0;
        end else begin
          regs_137_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_138_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h8a == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_138_0 <= 73'h0;
        end else begin
          regs_138_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_139_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h8b == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_139_0 <= 73'h0;
        end else begin
          regs_139_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_140_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h8c == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_140_0 <= 73'h0;
        end else begin
          regs_140_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_141_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h8d == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_141_0 <= 73'h0;
        end else begin
          regs_141_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_142_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h8e == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_142_0 <= 73'h0;
        end else begin
          regs_142_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_143_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h8f == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_143_0 <= 73'h0;
        end else begin
          regs_143_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_144_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h90 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_144_0 <= 73'h0;
        end else begin
          regs_144_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_145_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h91 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_145_0 <= 73'h0;
        end else begin
          regs_145_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_146_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h92 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_146_0 <= 73'h0;
        end else begin
          regs_146_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_147_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h93 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_147_0 <= 73'h0;
        end else begin
          regs_147_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_148_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h94 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_148_0 <= 73'h0;
        end else begin
          regs_148_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_149_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h95 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_149_0 <= 73'h0;
        end else begin
          regs_149_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_150_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h96 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_150_0 <= 73'h0;
        end else begin
          regs_150_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_151_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h97 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_151_0 <= 73'h0;
        end else begin
          regs_151_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_152_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h98 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_152_0 <= 73'h0;
        end else begin
          regs_152_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_153_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h99 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_153_0 <= 73'h0;
        end else begin
          regs_153_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_154_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h9a == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_154_0 <= 73'h0;
        end else begin
          regs_154_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_155_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h9b == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_155_0 <= 73'h0;
        end else begin
          regs_155_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_156_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h9c == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_156_0 <= 73'h0;
        end else begin
          regs_156_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_157_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h9d == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_157_0 <= 73'h0;
        end else begin
          regs_157_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_158_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h9e == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_158_0 <= 73'h0;
        end else begin
          regs_158_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_159_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h9f == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_159_0 <= 73'h0;
        end else begin
          regs_159_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_160_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'ha0 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_160_0 <= 73'h0;
        end else begin
          regs_160_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_161_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'ha1 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_161_0 <= 73'h0;
        end else begin
          regs_161_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_162_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'ha2 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_162_0 <= 73'h0;
        end else begin
          regs_162_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_163_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'ha3 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_163_0 <= 73'h0;
        end else begin
          regs_163_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_164_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'ha4 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_164_0 <= 73'h0;
        end else begin
          regs_164_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_165_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'ha5 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_165_0 <= 73'h0;
        end else begin
          regs_165_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_166_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'ha6 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_166_0 <= 73'h0;
        end else begin
          regs_166_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_167_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'ha7 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_167_0 <= 73'h0;
        end else begin
          regs_167_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_168_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'ha8 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_168_0 <= 73'h0;
        end else begin
          regs_168_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_169_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'ha9 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_169_0 <= 73'h0;
        end else begin
          regs_169_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_170_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'haa == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_170_0 <= 73'h0;
        end else begin
          regs_170_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_171_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hab == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_171_0 <= 73'h0;
        end else begin
          regs_171_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_172_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hac == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_172_0 <= 73'h0;
        end else begin
          regs_172_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_173_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'had == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_173_0 <= 73'h0;
        end else begin
          regs_173_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_174_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hae == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_174_0 <= 73'h0;
        end else begin
          regs_174_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_175_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'haf == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_175_0 <= 73'h0;
        end else begin
          regs_175_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_176_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hb0 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_176_0 <= 73'h0;
        end else begin
          regs_176_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_177_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hb1 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_177_0 <= 73'h0;
        end else begin
          regs_177_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_178_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hb2 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_178_0 <= 73'h0;
        end else begin
          regs_178_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_179_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hb3 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_179_0 <= 73'h0;
        end else begin
          regs_179_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_180_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hb4 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_180_0 <= 73'h0;
        end else begin
          regs_180_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_181_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hb5 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_181_0 <= 73'h0;
        end else begin
          regs_181_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_182_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hb6 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_182_0 <= 73'h0;
        end else begin
          regs_182_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_183_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hb7 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_183_0 <= 73'h0;
        end else begin
          regs_183_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_184_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hb8 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_184_0 <= 73'h0;
        end else begin
          regs_184_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_185_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hb9 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_185_0 <= 73'h0;
        end else begin
          regs_185_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_186_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hba == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_186_0 <= 73'h0;
        end else begin
          regs_186_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_187_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hbb == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_187_0 <= 73'h0;
        end else begin
          regs_187_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_188_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hbc == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_188_0 <= 73'h0;
        end else begin
          regs_188_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_189_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hbd == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_189_0 <= 73'h0;
        end else begin
          regs_189_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_190_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hbe == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_190_0 <= 73'h0;
        end else begin
          regs_190_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_191_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hbf == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_191_0 <= 73'h0;
        end else begin
          regs_191_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_192_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hc0 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_192_0 <= 73'h0;
        end else begin
          regs_192_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_193_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hc1 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_193_0 <= 73'h0;
        end else begin
          regs_193_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_194_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hc2 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_194_0 <= 73'h0;
        end else begin
          regs_194_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_195_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hc3 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_195_0 <= 73'h0;
        end else begin
          regs_195_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_196_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hc4 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_196_0 <= 73'h0;
        end else begin
          regs_196_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_197_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hc5 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_197_0 <= 73'h0;
        end else begin
          regs_197_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_198_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hc6 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_198_0 <= 73'h0;
        end else begin
          regs_198_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_199_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hc7 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_199_0 <= 73'h0;
        end else begin
          regs_199_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_200_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hc8 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_200_0 <= 73'h0;
        end else begin
          regs_200_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_201_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hc9 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_201_0 <= 73'h0;
        end else begin
          regs_201_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_202_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hca == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_202_0 <= 73'h0;
        end else begin
          regs_202_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_203_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hcb == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_203_0 <= 73'h0;
        end else begin
          regs_203_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_204_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hcc == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_204_0 <= 73'h0;
        end else begin
          regs_204_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_205_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hcd == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_205_0 <= 73'h0;
        end else begin
          regs_205_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_206_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hce == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_206_0 <= 73'h0;
        end else begin
          regs_206_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_207_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hcf == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_207_0 <= 73'h0;
        end else begin
          regs_207_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_208_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hd0 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_208_0 <= 73'h0;
        end else begin
          regs_208_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_209_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hd1 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_209_0 <= 73'h0;
        end else begin
          regs_209_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_210_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hd2 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_210_0 <= 73'h0;
        end else begin
          regs_210_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_211_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hd3 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_211_0 <= 73'h0;
        end else begin
          regs_211_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_212_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hd4 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_212_0 <= 73'h0;
        end else begin
          regs_212_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_213_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hd5 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_213_0 <= 73'h0;
        end else begin
          regs_213_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_214_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hd6 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_214_0 <= 73'h0;
        end else begin
          regs_214_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_215_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hd7 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_215_0 <= 73'h0;
        end else begin
          regs_215_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_216_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hd8 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_216_0 <= 73'h0;
        end else begin
          regs_216_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_217_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hd9 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_217_0 <= 73'h0;
        end else begin
          regs_217_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_218_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hda == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_218_0 <= 73'h0;
        end else begin
          regs_218_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_219_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hdb == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_219_0 <= 73'h0;
        end else begin
          regs_219_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_220_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hdc == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_220_0 <= 73'h0;
        end else begin
          regs_220_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_221_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hdd == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_221_0 <= 73'h0;
        end else begin
          regs_221_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_222_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hde == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_222_0 <= 73'h0;
        end else begin
          regs_222_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_223_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hdf == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_223_0 <= 73'h0;
        end else begin
          regs_223_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_224_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'he0 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_224_0 <= 73'h0;
        end else begin
          regs_224_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_225_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'he1 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_225_0 <= 73'h0;
        end else begin
          regs_225_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_226_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'he2 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_226_0 <= 73'h0;
        end else begin
          regs_226_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_227_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'he3 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_227_0 <= 73'h0;
        end else begin
          regs_227_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_228_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'he4 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_228_0 <= 73'h0;
        end else begin
          regs_228_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_229_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'he5 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_229_0 <= 73'h0;
        end else begin
          regs_229_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_230_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'he6 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_230_0 <= 73'h0;
        end else begin
          regs_230_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_231_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'he7 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_231_0 <= 73'h0;
        end else begin
          regs_231_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_232_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'he8 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_232_0 <= 73'h0;
        end else begin
          regs_232_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_233_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'he9 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_233_0 <= 73'h0;
        end else begin
          regs_233_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_234_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hea == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_234_0 <= 73'h0;
        end else begin
          regs_234_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_235_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'heb == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_235_0 <= 73'h0;
        end else begin
          regs_235_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_236_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hec == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_236_0 <= 73'h0;
        end else begin
          regs_236_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_237_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hed == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_237_0 <= 73'h0;
        end else begin
          regs_237_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_238_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hee == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_238_0 <= 73'h0;
        end else begin
          regs_238_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_239_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hef == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_239_0 <= 73'h0;
        end else begin
          regs_239_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_240_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hf0 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_240_0 <= 73'h0;
        end else begin
          regs_240_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_241_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hf1 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_241_0 <= 73'h0;
        end else begin
          regs_241_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_242_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hf2 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_242_0 <= 73'h0;
        end else begin
          regs_242_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_243_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hf3 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_243_0 <= 73'h0;
        end else begin
          regs_243_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_244_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hf4 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_244_0 <= 73'h0;
        end else begin
          regs_244_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_245_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hf5 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_245_0 <= 73'h0;
        end else begin
          regs_245_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_246_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hf6 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_246_0 <= 73'h0;
        end else begin
          regs_246_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_247_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hf7 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_247_0 <= 73'h0;
        end else begin
          regs_247_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_248_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hf8 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_248_0 <= 73'h0;
        end else begin
          regs_248_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_249_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hf9 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_249_0 <= 73'h0;
        end else begin
          regs_249_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_250_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hfa == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_250_0 <= 73'h0;
        end else begin
          regs_250_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_251_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hfb == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_251_0 <= 73'h0;
        end else begin
          regs_251_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_252_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hfc == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_252_0 <= 73'h0;
        end else begin
          regs_252_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_253_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hfd == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_253_0 <= 73'h0;
        end else begin
          regs_253_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_254_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hfe == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_254_0 <= 73'h0;
        end else begin
          regs_254_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_255_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'hff == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_255_0 <= 73'h0;
        end else begin
          regs_255_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_256_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h100 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_256_0 <= 73'h0;
        end else begin
          regs_256_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_257_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h101 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_257_0 <= 73'h0;
        end else begin
          regs_257_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_258_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h102 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_258_0 <= 73'h0;
        end else begin
          regs_258_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_259_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h103 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_259_0 <= 73'h0;
        end else begin
          regs_259_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_260_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h104 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_260_0 <= 73'h0;
        end else begin
          regs_260_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_261_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h105 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_261_0 <= 73'h0;
        end else begin
          regs_261_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_262_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h106 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_262_0 <= 73'h0;
        end else begin
          regs_262_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_263_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h107 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_263_0 <= 73'h0;
        end else begin
          regs_263_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_264_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h108 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_264_0 <= 73'h0;
        end else begin
          regs_264_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_265_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h109 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_265_0 <= 73'h0;
        end else begin
          regs_265_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_266_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h10a == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_266_0 <= 73'h0;
        end else begin
          regs_266_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_267_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h10b == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_267_0 <= 73'h0;
        end else begin
          regs_267_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_268_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h10c == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_268_0 <= 73'h0;
        end else begin
          regs_268_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_269_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h10d == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_269_0 <= 73'h0;
        end else begin
          regs_269_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_270_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h10e == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_270_0 <= 73'h0;
        end else begin
          regs_270_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_271_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h10f == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_271_0 <= 73'h0;
        end else begin
          regs_271_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_272_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h110 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_272_0 <= 73'h0;
        end else begin
          regs_272_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_273_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h111 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_273_0 <= 73'h0;
        end else begin
          regs_273_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_274_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h112 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_274_0 <= 73'h0;
        end else begin
          regs_274_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_275_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h113 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_275_0 <= 73'h0;
        end else begin
          regs_275_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_276_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h114 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_276_0 <= 73'h0;
        end else begin
          regs_276_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_277_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h115 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_277_0 <= 73'h0;
        end else begin
          regs_277_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_278_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h116 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_278_0 <= 73'h0;
        end else begin
          regs_278_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_279_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h117 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_279_0 <= 73'h0;
        end else begin
          regs_279_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_280_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h118 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_280_0 <= 73'h0;
        end else begin
          regs_280_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_281_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h119 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_281_0 <= 73'h0;
        end else begin
          regs_281_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_282_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h11a == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_282_0 <= 73'h0;
        end else begin
          regs_282_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_283_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h11b == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_283_0 <= 73'h0;
        end else begin
          regs_283_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_284_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h11c == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_284_0 <= 73'h0;
        end else begin
          regs_284_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_285_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h11d == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_285_0 <= 73'h0;
        end else begin
          regs_285_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_286_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h11e == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_286_0 <= 73'h0;
        end else begin
          regs_286_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_287_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h11f == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_287_0 <= 73'h0;
        end else begin
          regs_287_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_288_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h120 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_288_0 <= 73'h0;
        end else begin
          regs_288_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_289_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h121 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_289_0 <= 73'h0;
        end else begin
          regs_289_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_290_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h122 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_290_0 <= 73'h0;
        end else begin
          regs_290_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_291_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h123 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_291_0 <= 73'h0;
        end else begin
          regs_291_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_292_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h124 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_292_0 <= 73'h0;
        end else begin
          regs_292_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_293_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h125 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_293_0 <= 73'h0;
        end else begin
          regs_293_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_294_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h126 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_294_0 <= 73'h0;
        end else begin
          regs_294_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_295_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h127 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_295_0 <= 73'h0;
        end else begin
          regs_295_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_296_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h128 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_296_0 <= 73'h0;
        end else begin
          regs_296_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_297_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h129 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_297_0 <= 73'h0;
        end else begin
          regs_297_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_298_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h12a == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_298_0 <= 73'h0;
        end else begin
          regs_298_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_299_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h12b == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_299_0 <= 73'h0;
        end else begin
          regs_299_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_300_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h12c == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_300_0 <= 73'h0;
        end else begin
          regs_300_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_301_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h12d == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_301_0 <= 73'h0;
        end else begin
          regs_301_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_302_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h12e == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_302_0 <= 73'h0;
        end else begin
          regs_302_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_303_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h12f == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_303_0 <= 73'h0;
        end else begin
          regs_303_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_304_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h130 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_304_0 <= 73'h0;
        end else begin
          regs_304_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_305_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h131 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_305_0 <= 73'h0;
        end else begin
          regs_305_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_306_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h132 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_306_0 <= 73'h0;
        end else begin
          regs_306_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_307_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h133 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_307_0 <= 73'h0;
        end else begin
          regs_307_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_308_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h134 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_308_0 <= 73'h0;
        end else begin
          regs_308_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_309_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h135 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_309_0 <= 73'h0;
        end else begin
          regs_309_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_310_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h136 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_310_0 <= 73'h0;
        end else begin
          regs_310_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_311_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h137 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_311_0 <= 73'h0;
        end else begin
          regs_311_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_312_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h138 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_312_0 <= 73'h0;
        end else begin
          regs_312_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_313_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h139 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_313_0 <= 73'h0;
        end else begin
          regs_313_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_314_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h13a == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_314_0 <= 73'h0;
        end else begin
          regs_314_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_315_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h13b == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_315_0 <= 73'h0;
        end else begin
          regs_315_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_316_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h13c == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_316_0 <= 73'h0;
        end else begin
          regs_316_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_317_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h13d == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_317_0 <= 73'h0;
        end else begin
          regs_317_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_318_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h13e == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_318_0 <= 73'h0;
        end else begin
          regs_318_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_319_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h13f == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_319_0 <= 73'h0;
        end else begin
          regs_319_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_320_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h140 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_320_0 <= 73'h0;
        end else begin
          regs_320_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_321_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h141 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_321_0 <= 73'h0;
        end else begin
          regs_321_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_322_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h142 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_322_0 <= 73'h0;
        end else begin
          regs_322_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_323_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h143 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_323_0 <= 73'h0;
        end else begin
          regs_323_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_324_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h144 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_324_0 <= 73'h0;
        end else begin
          regs_324_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_325_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h145 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_325_0 <= 73'h0;
        end else begin
          regs_325_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_326_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h146 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_326_0 <= 73'h0;
        end else begin
          regs_326_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_327_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h147 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_327_0 <= 73'h0;
        end else begin
          regs_327_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_328_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h148 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_328_0 <= 73'h0;
        end else begin
          regs_328_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_329_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h149 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_329_0 <= 73'h0;
        end else begin
          regs_329_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_330_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h14a == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_330_0 <= 73'h0;
        end else begin
          regs_330_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_331_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h14b == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_331_0 <= 73'h0;
        end else begin
          regs_331_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_332_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h14c == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_332_0 <= 73'h0;
        end else begin
          regs_332_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_333_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h14d == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_333_0 <= 73'h0;
        end else begin
          regs_333_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_334_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h14e == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_334_0 <= 73'h0;
        end else begin
          regs_334_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_335_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h14f == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_335_0 <= 73'h0;
        end else begin
          regs_335_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_336_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h150 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_336_0 <= 73'h0;
        end else begin
          regs_336_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_337_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h151 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_337_0 <= 73'h0;
        end else begin
          regs_337_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_338_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h152 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_338_0 <= 73'h0;
        end else begin
          regs_338_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_339_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h153 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_339_0 <= 73'h0;
        end else begin
          regs_339_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_340_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h154 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_340_0 <= 73'h0;
        end else begin
          regs_340_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_341_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h155 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_341_0 <= 73'h0;
        end else begin
          regs_341_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_342_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h156 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_342_0 <= 73'h0;
        end else begin
          regs_342_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_343_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h157 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_343_0 <= 73'h0;
        end else begin
          regs_343_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_344_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h158 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_344_0 <= 73'h0;
        end else begin
          regs_344_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_345_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h159 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_345_0 <= 73'h0;
        end else begin
          regs_345_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_346_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h15a == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_346_0 <= 73'h0;
        end else begin
          regs_346_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_347_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h15b == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_347_0 <= 73'h0;
        end else begin
          regs_347_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_348_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h15c == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_348_0 <= 73'h0;
        end else begin
          regs_348_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_349_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h15d == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_349_0 <= 73'h0;
        end else begin
          regs_349_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_350_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h15e == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_350_0 <= 73'h0;
        end else begin
          regs_350_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_351_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h15f == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_351_0 <= 73'h0;
        end else begin
          regs_351_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_352_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h160 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_352_0 <= 73'h0;
        end else begin
          regs_352_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_353_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h161 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_353_0 <= 73'h0;
        end else begin
          regs_353_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_354_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h162 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_354_0 <= 73'h0;
        end else begin
          regs_354_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_355_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h163 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_355_0 <= 73'h0;
        end else begin
          regs_355_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_356_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h164 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_356_0 <= 73'h0;
        end else begin
          regs_356_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_357_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h165 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_357_0 <= 73'h0;
        end else begin
          regs_357_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_358_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h166 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_358_0 <= 73'h0;
        end else begin
          regs_358_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_359_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h167 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_359_0 <= 73'h0;
        end else begin
          regs_359_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_360_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h168 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_360_0 <= 73'h0;
        end else begin
          regs_360_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_361_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h169 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_361_0 <= 73'h0;
        end else begin
          regs_361_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_362_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h16a == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_362_0 <= 73'h0;
        end else begin
          regs_362_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_363_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h16b == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_363_0 <= 73'h0;
        end else begin
          regs_363_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_364_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h16c == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_364_0 <= 73'h0;
        end else begin
          regs_364_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_365_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h16d == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_365_0 <= 73'h0;
        end else begin
          regs_365_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_366_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h16e == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_366_0 <= 73'h0;
        end else begin
          regs_366_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_367_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h16f == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_367_0 <= 73'h0;
        end else begin
          regs_367_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_368_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h170 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_368_0 <= 73'h0;
        end else begin
          regs_368_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_369_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h171 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_369_0 <= 73'h0;
        end else begin
          regs_369_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_370_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h172 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_370_0 <= 73'h0;
        end else begin
          regs_370_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_371_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h173 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_371_0 <= 73'h0;
        end else begin
          regs_371_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_372_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h174 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_372_0 <= 73'h0;
        end else begin
          regs_372_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_373_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h175 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_373_0 <= 73'h0;
        end else begin
          regs_373_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_374_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h176 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_374_0 <= 73'h0;
        end else begin
          regs_374_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_375_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h177 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_375_0 <= 73'h0;
        end else begin
          regs_375_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_376_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h178 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_376_0 <= 73'h0;
        end else begin
          regs_376_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_377_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h179 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_377_0 <= 73'h0;
        end else begin
          regs_377_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_378_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h17a == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_378_0 <= 73'h0;
        end else begin
          regs_378_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_379_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h17b == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_379_0 <= 73'h0;
        end else begin
          regs_379_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_380_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h17c == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_380_0 <= 73'h0;
        end else begin
          regs_380_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_381_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h17d == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_381_0 <= 73'h0;
        end else begin
          regs_381_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_382_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h17e == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_382_0 <= 73'h0;
        end else begin
          regs_382_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_383_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h17f == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_383_0 <= 73'h0;
        end else begin
          regs_383_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_384_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h180 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_384_0 <= 73'h0;
        end else begin
          regs_384_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_385_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h181 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_385_0 <= 73'h0;
        end else begin
          regs_385_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_386_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h182 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_386_0 <= 73'h0;
        end else begin
          regs_386_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_387_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h183 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_387_0 <= 73'h0;
        end else begin
          regs_387_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_388_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h184 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_388_0 <= 73'h0;
        end else begin
          regs_388_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_389_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h185 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_389_0 <= 73'h0;
        end else begin
          regs_389_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_390_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h186 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_390_0 <= 73'h0;
        end else begin
          regs_390_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_391_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h187 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_391_0 <= 73'h0;
        end else begin
          regs_391_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_392_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h188 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_392_0 <= 73'h0;
        end else begin
          regs_392_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_393_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h189 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_393_0 <= 73'h0;
        end else begin
          regs_393_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_394_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h18a == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_394_0 <= 73'h0;
        end else begin
          regs_394_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_395_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h18b == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_395_0 <= 73'h0;
        end else begin
          regs_395_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_396_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h18c == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_396_0 <= 73'h0;
        end else begin
          regs_396_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_397_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h18d == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_397_0 <= 73'h0;
        end else begin
          regs_397_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_398_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h18e == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_398_0 <= 73'h0;
        end else begin
          regs_398_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_399_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h18f == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_399_0 <= 73'h0;
        end else begin
          regs_399_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_400_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h190 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_400_0 <= 73'h0;
        end else begin
          regs_400_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_401_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h191 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_401_0 <= 73'h0;
        end else begin
          regs_401_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_402_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h192 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_402_0 <= 73'h0;
        end else begin
          regs_402_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_403_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h193 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_403_0 <= 73'h0;
        end else begin
          regs_403_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_404_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h194 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_404_0 <= 73'h0;
        end else begin
          regs_404_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_405_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h195 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_405_0 <= 73'h0;
        end else begin
          regs_405_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_406_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h196 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_406_0 <= 73'h0;
        end else begin
          regs_406_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_407_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h197 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_407_0 <= 73'h0;
        end else begin
          regs_407_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_408_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h198 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_408_0 <= 73'h0;
        end else begin
          regs_408_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_409_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h199 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_409_0 <= 73'h0;
        end else begin
          regs_409_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_410_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h19a == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_410_0 <= 73'h0;
        end else begin
          regs_410_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_411_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h19b == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_411_0 <= 73'h0;
        end else begin
          regs_411_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_412_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h19c == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_412_0 <= 73'h0;
        end else begin
          regs_412_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_413_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h19d == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_413_0 <= 73'h0;
        end else begin
          regs_413_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_414_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h19e == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_414_0 <= 73'h0;
        end else begin
          regs_414_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_415_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h19f == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_415_0 <= 73'h0;
        end else begin
          regs_415_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_416_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1a0 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_416_0 <= 73'h0;
        end else begin
          regs_416_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_417_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1a1 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_417_0 <= 73'h0;
        end else begin
          regs_417_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_418_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1a2 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_418_0 <= 73'h0;
        end else begin
          regs_418_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_419_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1a3 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_419_0 <= 73'h0;
        end else begin
          regs_419_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_420_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1a4 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_420_0 <= 73'h0;
        end else begin
          regs_420_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_421_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1a5 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_421_0 <= 73'h0;
        end else begin
          regs_421_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_422_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1a6 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_422_0 <= 73'h0;
        end else begin
          regs_422_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_423_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1a7 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_423_0 <= 73'h0;
        end else begin
          regs_423_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_424_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1a8 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_424_0 <= 73'h0;
        end else begin
          regs_424_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_425_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1a9 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_425_0 <= 73'h0;
        end else begin
          regs_425_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_426_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1aa == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_426_0 <= 73'h0;
        end else begin
          regs_426_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_427_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1ab == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_427_0 <= 73'h0;
        end else begin
          regs_427_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_428_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1ac == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_428_0 <= 73'h0;
        end else begin
          regs_428_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_429_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1ad == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_429_0 <= 73'h0;
        end else begin
          regs_429_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_430_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1ae == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_430_0 <= 73'h0;
        end else begin
          regs_430_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_431_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1af == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_431_0 <= 73'h0;
        end else begin
          regs_431_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_432_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1b0 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_432_0 <= 73'h0;
        end else begin
          regs_432_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_433_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1b1 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_433_0 <= 73'h0;
        end else begin
          regs_433_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_434_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1b2 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_434_0 <= 73'h0;
        end else begin
          regs_434_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_435_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1b3 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_435_0 <= 73'h0;
        end else begin
          regs_435_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_436_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1b4 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_436_0 <= 73'h0;
        end else begin
          regs_436_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_437_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1b5 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_437_0 <= 73'h0;
        end else begin
          regs_437_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_438_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1b6 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_438_0 <= 73'h0;
        end else begin
          regs_438_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_439_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1b7 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_439_0 <= 73'h0;
        end else begin
          regs_439_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_440_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1b8 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_440_0 <= 73'h0;
        end else begin
          regs_440_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_441_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1b9 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_441_0 <= 73'h0;
        end else begin
          regs_441_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_442_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1ba == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_442_0 <= 73'h0;
        end else begin
          regs_442_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_443_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1bb == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_443_0 <= 73'h0;
        end else begin
          regs_443_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_444_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1bc == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_444_0 <= 73'h0;
        end else begin
          regs_444_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_445_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1bd == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_445_0 <= 73'h0;
        end else begin
          regs_445_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_446_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1be == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_446_0 <= 73'h0;
        end else begin
          regs_446_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_447_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1bf == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_447_0 <= 73'h0;
        end else begin
          regs_447_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_448_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1c0 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_448_0 <= 73'h0;
        end else begin
          regs_448_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_449_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1c1 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_449_0 <= 73'h0;
        end else begin
          regs_449_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_450_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1c2 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_450_0 <= 73'h0;
        end else begin
          regs_450_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_451_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1c3 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_451_0 <= 73'h0;
        end else begin
          regs_451_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_452_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1c4 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_452_0 <= 73'h0;
        end else begin
          regs_452_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_453_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1c5 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_453_0 <= 73'h0;
        end else begin
          regs_453_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_454_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1c6 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_454_0 <= 73'h0;
        end else begin
          regs_454_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_455_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1c7 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_455_0 <= 73'h0;
        end else begin
          regs_455_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_456_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1c8 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_456_0 <= 73'h0;
        end else begin
          regs_456_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_457_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1c9 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_457_0 <= 73'h0;
        end else begin
          regs_457_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_458_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1ca == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_458_0 <= 73'h0;
        end else begin
          regs_458_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_459_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1cb == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_459_0 <= 73'h0;
        end else begin
          regs_459_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_460_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1cc == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_460_0 <= 73'h0;
        end else begin
          regs_460_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_461_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1cd == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_461_0 <= 73'h0;
        end else begin
          regs_461_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_462_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1ce == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_462_0 <= 73'h0;
        end else begin
          regs_462_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_463_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1cf == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_463_0 <= 73'h0;
        end else begin
          regs_463_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_464_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1d0 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_464_0 <= 73'h0;
        end else begin
          regs_464_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_465_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1d1 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_465_0 <= 73'h0;
        end else begin
          regs_465_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_466_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1d2 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_466_0 <= 73'h0;
        end else begin
          regs_466_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_467_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1d3 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_467_0 <= 73'h0;
        end else begin
          regs_467_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_468_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1d4 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_468_0 <= 73'h0;
        end else begin
          regs_468_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_469_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1d5 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_469_0 <= 73'h0;
        end else begin
          regs_469_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_470_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1d6 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_470_0 <= 73'h0;
        end else begin
          regs_470_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_471_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1d7 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_471_0 <= 73'h0;
        end else begin
          regs_471_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_472_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1d8 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_472_0 <= 73'h0;
        end else begin
          regs_472_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_473_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1d9 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_473_0 <= 73'h0;
        end else begin
          regs_473_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_474_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1da == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_474_0 <= 73'h0;
        end else begin
          regs_474_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_475_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1db == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_475_0 <= 73'h0;
        end else begin
          regs_475_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_476_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1dc == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_476_0 <= 73'h0;
        end else begin
          regs_476_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_477_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1dd == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_477_0 <= 73'h0;
        end else begin
          regs_477_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_478_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1de == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_478_0 <= 73'h0;
        end else begin
          regs_478_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_479_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1df == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_479_0 <= 73'h0;
        end else begin
          regs_479_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_480_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1e0 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_480_0 <= 73'h0;
        end else begin
          regs_480_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_481_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1e1 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_481_0 <= 73'h0;
        end else begin
          regs_481_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_482_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1e2 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_482_0 <= 73'h0;
        end else begin
          regs_482_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_483_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1e3 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_483_0 <= 73'h0;
        end else begin
          regs_483_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_484_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1e4 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_484_0 <= 73'h0;
        end else begin
          regs_484_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_485_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1e5 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_485_0 <= 73'h0;
        end else begin
          regs_485_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_486_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1e6 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_486_0 <= 73'h0;
        end else begin
          regs_486_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_487_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1e7 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_487_0 <= 73'h0;
        end else begin
          regs_487_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_488_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1e8 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_488_0 <= 73'h0;
        end else begin
          regs_488_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_489_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1e9 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_489_0 <= 73'h0;
        end else begin
          regs_489_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_490_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1ea == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_490_0 <= 73'h0;
        end else begin
          regs_490_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_491_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1eb == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_491_0 <= 73'h0;
        end else begin
          regs_491_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_492_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1ec == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_492_0 <= 73'h0;
        end else begin
          regs_492_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_493_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1ed == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_493_0 <= 73'h0;
        end else begin
          regs_493_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_494_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1ee == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_494_0 <= 73'h0;
        end else begin
          regs_494_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_495_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1ef == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_495_0 <= 73'h0;
        end else begin
          regs_495_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_496_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1f0 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_496_0 <= 73'h0;
        end else begin
          regs_496_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_497_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1f1 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_497_0 <= 73'h0;
        end else begin
          regs_497_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_498_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1f2 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_498_0 <= 73'h0;
        end else begin
          regs_498_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_499_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1f3 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_499_0 <= 73'h0;
        end else begin
          regs_499_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_500_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1f4 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_500_0 <= 73'h0;
        end else begin
          regs_500_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_501_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1f5 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_501_0 <= 73'h0;
        end else begin
          regs_501_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_502_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1f6 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_502_0 <= 73'h0;
        end else begin
          regs_502_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_503_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1f7 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_503_0 <= 73'h0;
        end else begin
          regs_503_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_504_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1f8 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_504_0 <= 73'h0;
        end else begin
          regs_504_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_505_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1f9 == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_505_0 <= 73'h0;
        end else begin
          regs_505_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_506_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1fa == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_506_0 <= 73'h0;
        end else begin
          regs_506_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_507_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1fb == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_507_0 <= 73'h0;
        end else begin
          regs_507_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_508_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1fc == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_508_0 <= 73'h0;
        end else begin
          regs_508_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_509_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1fd == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_509_0 <= 73'h0;
        end else begin
          regs_509_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_510_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1fe == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_510_0 <= 73'h0;
        end else begin
          regs_510_0 <= _wdataword_T;
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_511_0 <= 73'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (wen) begin // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
      if (9'h1ff == setIdx) begin // @[src/main/scala/utils/RegMem.scala 22:21]
        if (resetState) begin // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
          regs_511_0 <= 73'h0;
        end else begin
          regs_511_0 <= _wdataword_T;
        end
      end
    end
    resetState <= reset | _GEN_2; // @[src/main/scala/utils/SRAMTemplate.scala 80:{30,30}]
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      resetSet <= 9'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (resetState) begin // @[src/main/scala/chisel3/util/Counter.scala 118:16]
      resetSet <= _wrap_value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (realRen) begin // @[src/main/scala/utils/RegMem.scala 39:14]
      if (9'h1ff == io_r_req_bits_setIdx) begin // @[src/main/scala/utils/RegMem.scala 39:14]
        rdata_r_0 <= regs_511_0; // @[src/main/scala/utils/RegMem.scala 39:14]
      end else if (9'h1fe == io_r_req_bits_setIdx) begin // @[src/main/scala/utils/RegMem.scala 39:14]
        rdata_r_0 <= regs_510_0; // @[src/main/scala/utils/RegMem.scala 39:14]
      end else if (9'h1fd == io_r_req_bits_setIdx) begin // @[src/main/scala/utils/RegMem.scala 39:14]
        rdata_r_0 <= regs_509_0; // @[src/main/scala/utils/RegMem.scala 39:14]
      end else begin
        rdata_r_0 <= _GEN_2047;
      end
    end
    rdata_REG <= io_r_req_valid & ~wen; // @[src/main/scala/utils/SRAMTemplate.scala 89:38]
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      rdata_r_1_0 <= 73'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (rdata_REG) begin // @[src/main/scala/utils/Hold.scala 23:65]
      rdata_r_1_0 <= rdata_r_0; // @[src/main/scala/utils/Hold.scala 23:65]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {3{`RANDOM}};
  regs_0_0 = _RAND_0[72:0];
  _RAND_1 = {3{`RANDOM}};
  regs_1_0 = _RAND_1[72:0];
  _RAND_2 = {3{`RANDOM}};
  regs_2_0 = _RAND_2[72:0];
  _RAND_3 = {3{`RANDOM}};
  regs_3_0 = _RAND_3[72:0];
  _RAND_4 = {3{`RANDOM}};
  regs_4_0 = _RAND_4[72:0];
  _RAND_5 = {3{`RANDOM}};
  regs_5_0 = _RAND_5[72:0];
  _RAND_6 = {3{`RANDOM}};
  regs_6_0 = _RAND_6[72:0];
  _RAND_7 = {3{`RANDOM}};
  regs_7_0 = _RAND_7[72:0];
  _RAND_8 = {3{`RANDOM}};
  regs_8_0 = _RAND_8[72:0];
  _RAND_9 = {3{`RANDOM}};
  regs_9_0 = _RAND_9[72:0];
  _RAND_10 = {3{`RANDOM}};
  regs_10_0 = _RAND_10[72:0];
  _RAND_11 = {3{`RANDOM}};
  regs_11_0 = _RAND_11[72:0];
  _RAND_12 = {3{`RANDOM}};
  regs_12_0 = _RAND_12[72:0];
  _RAND_13 = {3{`RANDOM}};
  regs_13_0 = _RAND_13[72:0];
  _RAND_14 = {3{`RANDOM}};
  regs_14_0 = _RAND_14[72:0];
  _RAND_15 = {3{`RANDOM}};
  regs_15_0 = _RAND_15[72:0];
  _RAND_16 = {3{`RANDOM}};
  regs_16_0 = _RAND_16[72:0];
  _RAND_17 = {3{`RANDOM}};
  regs_17_0 = _RAND_17[72:0];
  _RAND_18 = {3{`RANDOM}};
  regs_18_0 = _RAND_18[72:0];
  _RAND_19 = {3{`RANDOM}};
  regs_19_0 = _RAND_19[72:0];
  _RAND_20 = {3{`RANDOM}};
  regs_20_0 = _RAND_20[72:0];
  _RAND_21 = {3{`RANDOM}};
  regs_21_0 = _RAND_21[72:0];
  _RAND_22 = {3{`RANDOM}};
  regs_22_0 = _RAND_22[72:0];
  _RAND_23 = {3{`RANDOM}};
  regs_23_0 = _RAND_23[72:0];
  _RAND_24 = {3{`RANDOM}};
  regs_24_0 = _RAND_24[72:0];
  _RAND_25 = {3{`RANDOM}};
  regs_25_0 = _RAND_25[72:0];
  _RAND_26 = {3{`RANDOM}};
  regs_26_0 = _RAND_26[72:0];
  _RAND_27 = {3{`RANDOM}};
  regs_27_0 = _RAND_27[72:0];
  _RAND_28 = {3{`RANDOM}};
  regs_28_0 = _RAND_28[72:0];
  _RAND_29 = {3{`RANDOM}};
  regs_29_0 = _RAND_29[72:0];
  _RAND_30 = {3{`RANDOM}};
  regs_30_0 = _RAND_30[72:0];
  _RAND_31 = {3{`RANDOM}};
  regs_31_0 = _RAND_31[72:0];
  _RAND_32 = {3{`RANDOM}};
  regs_32_0 = _RAND_32[72:0];
  _RAND_33 = {3{`RANDOM}};
  regs_33_0 = _RAND_33[72:0];
  _RAND_34 = {3{`RANDOM}};
  regs_34_0 = _RAND_34[72:0];
  _RAND_35 = {3{`RANDOM}};
  regs_35_0 = _RAND_35[72:0];
  _RAND_36 = {3{`RANDOM}};
  regs_36_0 = _RAND_36[72:0];
  _RAND_37 = {3{`RANDOM}};
  regs_37_0 = _RAND_37[72:0];
  _RAND_38 = {3{`RANDOM}};
  regs_38_0 = _RAND_38[72:0];
  _RAND_39 = {3{`RANDOM}};
  regs_39_0 = _RAND_39[72:0];
  _RAND_40 = {3{`RANDOM}};
  regs_40_0 = _RAND_40[72:0];
  _RAND_41 = {3{`RANDOM}};
  regs_41_0 = _RAND_41[72:0];
  _RAND_42 = {3{`RANDOM}};
  regs_42_0 = _RAND_42[72:0];
  _RAND_43 = {3{`RANDOM}};
  regs_43_0 = _RAND_43[72:0];
  _RAND_44 = {3{`RANDOM}};
  regs_44_0 = _RAND_44[72:0];
  _RAND_45 = {3{`RANDOM}};
  regs_45_0 = _RAND_45[72:0];
  _RAND_46 = {3{`RANDOM}};
  regs_46_0 = _RAND_46[72:0];
  _RAND_47 = {3{`RANDOM}};
  regs_47_0 = _RAND_47[72:0];
  _RAND_48 = {3{`RANDOM}};
  regs_48_0 = _RAND_48[72:0];
  _RAND_49 = {3{`RANDOM}};
  regs_49_0 = _RAND_49[72:0];
  _RAND_50 = {3{`RANDOM}};
  regs_50_0 = _RAND_50[72:0];
  _RAND_51 = {3{`RANDOM}};
  regs_51_0 = _RAND_51[72:0];
  _RAND_52 = {3{`RANDOM}};
  regs_52_0 = _RAND_52[72:0];
  _RAND_53 = {3{`RANDOM}};
  regs_53_0 = _RAND_53[72:0];
  _RAND_54 = {3{`RANDOM}};
  regs_54_0 = _RAND_54[72:0];
  _RAND_55 = {3{`RANDOM}};
  regs_55_0 = _RAND_55[72:0];
  _RAND_56 = {3{`RANDOM}};
  regs_56_0 = _RAND_56[72:0];
  _RAND_57 = {3{`RANDOM}};
  regs_57_0 = _RAND_57[72:0];
  _RAND_58 = {3{`RANDOM}};
  regs_58_0 = _RAND_58[72:0];
  _RAND_59 = {3{`RANDOM}};
  regs_59_0 = _RAND_59[72:0];
  _RAND_60 = {3{`RANDOM}};
  regs_60_0 = _RAND_60[72:0];
  _RAND_61 = {3{`RANDOM}};
  regs_61_0 = _RAND_61[72:0];
  _RAND_62 = {3{`RANDOM}};
  regs_62_0 = _RAND_62[72:0];
  _RAND_63 = {3{`RANDOM}};
  regs_63_0 = _RAND_63[72:0];
  _RAND_64 = {3{`RANDOM}};
  regs_64_0 = _RAND_64[72:0];
  _RAND_65 = {3{`RANDOM}};
  regs_65_0 = _RAND_65[72:0];
  _RAND_66 = {3{`RANDOM}};
  regs_66_0 = _RAND_66[72:0];
  _RAND_67 = {3{`RANDOM}};
  regs_67_0 = _RAND_67[72:0];
  _RAND_68 = {3{`RANDOM}};
  regs_68_0 = _RAND_68[72:0];
  _RAND_69 = {3{`RANDOM}};
  regs_69_0 = _RAND_69[72:0];
  _RAND_70 = {3{`RANDOM}};
  regs_70_0 = _RAND_70[72:0];
  _RAND_71 = {3{`RANDOM}};
  regs_71_0 = _RAND_71[72:0];
  _RAND_72 = {3{`RANDOM}};
  regs_72_0 = _RAND_72[72:0];
  _RAND_73 = {3{`RANDOM}};
  regs_73_0 = _RAND_73[72:0];
  _RAND_74 = {3{`RANDOM}};
  regs_74_0 = _RAND_74[72:0];
  _RAND_75 = {3{`RANDOM}};
  regs_75_0 = _RAND_75[72:0];
  _RAND_76 = {3{`RANDOM}};
  regs_76_0 = _RAND_76[72:0];
  _RAND_77 = {3{`RANDOM}};
  regs_77_0 = _RAND_77[72:0];
  _RAND_78 = {3{`RANDOM}};
  regs_78_0 = _RAND_78[72:0];
  _RAND_79 = {3{`RANDOM}};
  regs_79_0 = _RAND_79[72:0];
  _RAND_80 = {3{`RANDOM}};
  regs_80_0 = _RAND_80[72:0];
  _RAND_81 = {3{`RANDOM}};
  regs_81_0 = _RAND_81[72:0];
  _RAND_82 = {3{`RANDOM}};
  regs_82_0 = _RAND_82[72:0];
  _RAND_83 = {3{`RANDOM}};
  regs_83_0 = _RAND_83[72:0];
  _RAND_84 = {3{`RANDOM}};
  regs_84_0 = _RAND_84[72:0];
  _RAND_85 = {3{`RANDOM}};
  regs_85_0 = _RAND_85[72:0];
  _RAND_86 = {3{`RANDOM}};
  regs_86_0 = _RAND_86[72:0];
  _RAND_87 = {3{`RANDOM}};
  regs_87_0 = _RAND_87[72:0];
  _RAND_88 = {3{`RANDOM}};
  regs_88_0 = _RAND_88[72:0];
  _RAND_89 = {3{`RANDOM}};
  regs_89_0 = _RAND_89[72:0];
  _RAND_90 = {3{`RANDOM}};
  regs_90_0 = _RAND_90[72:0];
  _RAND_91 = {3{`RANDOM}};
  regs_91_0 = _RAND_91[72:0];
  _RAND_92 = {3{`RANDOM}};
  regs_92_0 = _RAND_92[72:0];
  _RAND_93 = {3{`RANDOM}};
  regs_93_0 = _RAND_93[72:0];
  _RAND_94 = {3{`RANDOM}};
  regs_94_0 = _RAND_94[72:0];
  _RAND_95 = {3{`RANDOM}};
  regs_95_0 = _RAND_95[72:0];
  _RAND_96 = {3{`RANDOM}};
  regs_96_0 = _RAND_96[72:0];
  _RAND_97 = {3{`RANDOM}};
  regs_97_0 = _RAND_97[72:0];
  _RAND_98 = {3{`RANDOM}};
  regs_98_0 = _RAND_98[72:0];
  _RAND_99 = {3{`RANDOM}};
  regs_99_0 = _RAND_99[72:0];
  _RAND_100 = {3{`RANDOM}};
  regs_100_0 = _RAND_100[72:0];
  _RAND_101 = {3{`RANDOM}};
  regs_101_0 = _RAND_101[72:0];
  _RAND_102 = {3{`RANDOM}};
  regs_102_0 = _RAND_102[72:0];
  _RAND_103 = {3{`RANDOM}};
  regs_103_0 = _RAND_103[72:0];
  _RAND_104 = {3{`RANDOM}};
  regs_104_0 = _RAND_104[72:0];
  _RAND_105 = {3{`RANDOM}};
  regs_105_0 = _RAND_105[72:0];
  _RAND_106 = {3{`RANDOM}};
  regs_106_0 = _RAND_106[72:0];
  _RAND_107 = {3{`RANDOM}};
  regs_107_0 = _RAND_107[72:0];
  _RAND_108 = {3{`RANDOM}};
  regs_108_0 = _RAND_108[72:0];
  _RAND_109 = {3{`RANDOM}};
  regs_109_0 = _RAND_109[72:0];
  _RAND_110 = {3{`RANDOM}};
  regs_110_0 = _RAND_110[72:0];
  _RAND_111 = {3{`RANDOM}};
  regs_111_0 = _RAND_111[72:0];
  _RAND_112 = {3{`RANDOM}};
  regs_112_0 = _RAND_112[72:0];
  _RAND_113 = {3{`RANDOM}};
  regs_113_0 = _RAND_113[72:0];
  _RAND_114 = {3{`RANDOM}};
  regs_114_0 = _RAND_114[72:0];
  _RAND_115 = {3{`RANDOM}};
  regs_115_0 = _RAND_115[72:0];
  _RAND_116 = {3{`RANDOM}};
  regs_116_0 = _RAND_116[72:0];
  _RAND_117 = {3{`RANDOM}};
  regs_117_0 = _RAND_117[72:0];
  _RAND_118 = {3{`RANDOM}};
  regs_118_0 = _RAND_118[72:0];
  _RAND_119 = {3{`RANDOM}};
  regs_119_0 = _RAND_119[72:0];
  _RAND_120 = {3{`RANDOM}};
  regs_120_0 = _RAND_120[72:0];
  _RAND_121 = {3{`RANDOM}};
  regs_121_0 = _RAND_121[72:0];
  _RAND_122 = {3{`RANDOM}};
  regs_122_0 = _RAND_122[72:0];
  _RAND_123 = {3{`RANDOM}};
  regs_123_0 = _RAND_123[72:0];
  _RAND_124 = {3{`RANDOM}};
  regs_124_0 = _RAND_124[72:0];
  _RAND_125 = {3{`RANDOM}};
  regs_125_0 = _RAND_125[72:0];
  _RAND_126 = {3{`RANDOM}};
  regs_126_0 = _RAND_126[72:0];
  _RAND_127 = {3{`RANDOM}};
  regs_127_0 = _RAND_127[72:0];
  _RAND_128 = {3{`RANDOM}};
  regs_128_0 = _RAND_128[72:0];
  _RAND_129 = {3{`RANDOM}};
  regs_129_0 = _RAND_129[72:0];
  _RAND_130 = {3{`RANDOM}};
  regs_130_0 = _RAND_130[72:0];
  _RAND_131 = {3{`RANDOM}};
  regs_131_0 = _RAND_131[72:0];
  _RAND_132 = {3{`RANDOM}};
  regs_132_0 = _RAND_132[72:0];
  _RAND_133 = {3{`RANDOM}};
  regs_133_0 = _RAND_133[72:0];
  _RAND_134 = {3{`RANDOM}};
  regs_134_0 = _RAND_134[72:0];
  _RAND_135 = {3{`RANDOM}};
  regs_135_0 = _RAND_135[72:0];
  _RAND_136 = {3{`RANDOM}};
  regs_136_0 = _RAND_136[72:0];
  _RAND_137 = {3{`RANDOM}};
  regs_137_0 = _RAND_137[72:0];
  _RAND_138 = {3{`RANDOM}};
  regs_138_0 = _RAND_138[72:0];
  _RAND_139 = {3{`RANDOM}};
  regs_139_0 = _RAND_139[72:0];
  _RAND_140 = {3{`RANDOM}};
  regs_140_0 = _RAND_140[72:0];
  _RAND_141 = {3{`RANDOM}};
  regs_141_0 = _RAND_141[72:0];
  _RAND_142 = {3{`RANDOM}};
  regs_142_0 = _RAND_142[72:0];
  _RAND_143 = {3{`RANDOM}};
  regs_143_0 = _RAND_143[72:0];
  _RAND_144 = {3{`RANDOM}};
  regs_144_0 = _RAND_144[72:0];
  _RAND_145 = {3{`RANDOM}};
  regs_145_0 = _RAND_145[72:0];
  _RAND_146 = {3{`RANDOM}};
  regs_146_0 = _RAND_146[72:0];
  _RAND_147 = {3{`RANDOM}};
  regs_147_0 = _RAND_147[72:0];
  _RAND_148 = {3{`RANDOM}};
  regs_148_0 = _RAND_148[72:0];
  _RAND_149 = {3{`RANDOM}};
  regs_149_0 = _RAND_149[72:0];
  _RAND_150 = {3{`RANDOM}};
  regs_150_0 = _RAND_150[72:0];
  _RAND_151 = {3{`RANDOM}};
  regs_151_0 = _RAND_151[72:0];
  _RAND_152 = {3{`RANDOM}};
  regs_152_0 = _RAND_152[72:0];
  _RAND_153 = {3{`RANDOM}};
  regs_153_0 = _RAND_153[72:0];
  _RAND_154 = {3{`RANDOM}};
  regs_154_0 = _RAND_154[72:0];
  _RAND_155 = {3{`RANDOM}};
  regs_155_0 = _RAND_155[72:0];
  _RAND_156 = {3{`RANDOM}};
  regs_156_0 = _RAND_156[72:0];
  _RAND_157 = {3{`RANDOM}};
  regs_157_0 = _RAND_157[72:0];
  _RAND_158 = {3{`RANDOM}};
  regs_158_0 = _RAND_158[72:0];
  _RAND_159 = {3{`RANDOM}};
  regs_159_0 = _RAND_159[72:0];
  _RAND_160 = {3{`RANDOM}};
  regs_160_0 = _RAND_160[72:0];
  _RAND_161 = {3{`RANDOM}};
  regs_161_0 = _RAND_161[72:0];
  _RAND_162 = {3{`RANDOM}};
  regs_162_0 = _RAND_162[72:0];
  _RAND_163 = {3{`RANDOM}};
  regs_163_0 = _RAND_163[72:0];
  _RAND_164 = {3{`RANDOM}};
  regs_164_0 = _RAND_164[72:0];
  _RAND_165 = {3{`RANDOM}};
  regs_165_0 = _RAND_165[72:0];
  _RAND_166 = {3{`RANDOM}};
  regs_166_0 = _RAND_166[72:0];
  _RAND_167 = {3{`RANDOM}};
  regs_167_0 = _RAND_167[72:0];
  _RAND_168 = {3{`RANDOM}};
  regs_168_0 = _RAND_168[72:0];
  _RAND_169 = {3{`RANDOM}};
  regs_169_0 = _RAND_169[72:0];
  _RAND_170 = {3{`RANDOM}};
  regs_170_0 = _RAND_170[72:0];
  _RAND_171 = {3{`RANDOM}};
  regs_171_0 = _RAND_171[72:0];
  _RAND_172 = {3{`RANDOM}};
  regs_172_0 = _RAND_172[72:0];
  _RAND_173 = {3{`RANDOM}};
  regs_173_0 = _RAND_173[72:0];
  _RAND_174 = {3{`RANDOM}};
  regs_174_0 = _RAND_174[72:0];
  _RAND_175 = {3{`RANDOM}};
  regs_175_0 = _RAND_175[72:0];
  _RAND_176 = {3{`RANDOM}};
  regs_176_0 = _RAND_176[72:0];
  _RAND_177 = {3{`RANDOM}};
  regs_177_0 = _RAND_177[72:0];
  _RAND_178 = {3{`RANDOM}};
  regs_178_0 = _RAND_178[72:0];
  _RAND_179 = {3{`RANDOM}};
  regs_179_0 = _RAND_179[72:0];
  _RAND_180 = {3{`RANDOM}};
  regs_180_0 = _RAND_180[72:0];
  _RAND_181 = {3{`RANDOM}};
  regs_181_0 = _RAND_181[72:0];
  _RAND_182 = {3{`RANDOM}};
  regs_182_0 = _RAND_182[72:0];
  _RAND_183 = {3{`RANDOM}};
  regs_183_0 = _RAND_183[72:0];
  _RAND_184 = {3{`RANDOM}};
  regs_184_0 = _RAND_184[72:0];
  _RAND_185 = {3{`RANDOM}};
  regs_185_0 = _RAND_185[72:0];
  _RAND_186 = {3{`RANDOM}};
  regs_186_0 = _RAND_186[72:0];
  _RAND_187 = {3{`RANDOM}};
  regs_187_0 = _RAND_187[72:0];
  _RAND_188 = {3{`RANDOM}};
  regs_188_0 = _RAND_188[72:0];
  _RAND_189 = {3{`RANDOM}};
  regs_189_0 = _RAND_189[72:0];
  _RAND_190 = {3{`RANDOM}};
  regs_190_0 = _RAND_190[72:0];
  _RAND_191 = {3{`RANDOM}};
  regs_191_0 = _RAND_191[72:0];
  _RAND_192 = {3{`RANDOM}};
  regs_192_0 = _RAND_192[72:0];
  _RAND_193 = {3{`RANDOM}};
  regs_193_0 = _RAND_193[72:0];
  _RAND_194 = {3{`RANDOM}};
  regs_194_0 = _RAND_194[72:0];
  _RAND_195 = {3{`RANDOM}};
  regs_195_0 = _RAND_195[72:0];
  _RAND_196 = {3{`RANDOM}};
  regs_196_0 = _RAND_196[72:0];
  _RAND_197 = {3{`RANDOM}};
  regs_197_0 = _RAND_197[72:0];
  _RAND_198 = {3{`RANDOM}};
  regs_198_0 = _RAND_198[72:0];
  _RAND_199 = {3{`RANDOM}};
  regs_199_0 = _RAND_199[72:0];
  _RAND_200 = {3{`RANDOM}};
  regs_200_0 = _RAND_200[72:0];
  _RAND_201 = {3{`RANDOM}};
  regs_201_0 = _RAND_201[72:0];
  _RAND_202 = {3{`RANDOM}};
  regs_202_0 = _RAND_202[72:0];
  _RAND_203 = {3{`RANDOM}};
  regs_203_0 = _RAND_203[72:0];
  _RAND_204 = {3{`RANDOM}};
  regs_204_0 = _RAND_204[72:0];
  _RAND_205 = {3{`RANDOM}};
  regs_205_0 = _RAND_205[72:0];
  _RAND_206 = {3{`RANDOM}};
  regs_206_0 = _RAND_206[72:0];
  _RAND_207 = {3{`RANDOM}};
  regs_207_0 = _RAND_207[72:0];
  _RAND_208 = {3{`RANDOM}};
  regs_208_0 = _RAND_208[72:0];
  _RAND_209 = {3{`RANDOM}};
  regs_209_0 = _RAND_209[72:0];
  _RAND_210 = {3{`RANDOM}};
  regs_210_0 = _RAND_210[72:0];
  _RAND_211 = {3{`RANDOM}};
  regs_211_0 = _RAND_211[72:0];
  _RAND_212 = {3{`RANDOM}};
  regs_212_0 = _RAND_212[72:0];
  _RAND_213 = {3{`RANDOM}};
  regs_213_0 = _RAND_213[72:0];
  _RAND_214 = {3{`RANDOM}};
  regs_214_0 = _RAND_214[72:0];
  _RAND_215 = {3{`RANDOM}};
  regs_215_0 = _RAND_215[72:0];
  _RAND_216 = {3{`RANDOM}};
  regs_216_0 = _RAND_216[72:0];
  _RAND_217 = {3{`RANDOM}};
  regs_217_0 = _RAND_217[72:0];
  _RAND_218 = {3{`RANDOM}};
  regs_218_0 = _RAND_218[72:0];
  _RAND_219 = {3{`RANDOM}};
  regs_219_0 = _RAND_219[72:0];
  _RAND_220 = {3{`RANDOM}};
  regs_220_0 = _RAND_220[72:0];
  _RAND_221 = {3{`RANDOM}};
  regs_221_0 = _RAND_221[72:0];
  _RAND_222 = {3{`RANDOM}};
  regs_222_0 = _RAND_222[72:0];
  _RAND_223 = {3{`RANDOM}};
  regs_223_0 = _RAND_223[72:0];
  _RAND_224 = {3{`RANDOM}};
  regs_224_0 = _RAND_224[72:0];
  _RAND_225 = {3{`RANDOM}};
  regs_225_0 = _RAND_225[72:0];
  _RAND_226 = {3{`RANDOM}};
  regs_226_0 = _RAND_226[72:0];
  _RAND_227 = {3{`RANDOM}};
  regs_227_0 = _RAND_227[72:0];
  _RAND_228 = {3{`RANDOM}};
  regs_228_0 = _RAND_228[72:0];
  _RAND_229 = {3{`RANDOM}};
  regs_229_0 = _RAND_229[72:0];
  _RAND_230 = {3{`RANDOM}};
  regs_230_0 = _RAND_230[72:0];
  _RAND_231 = {3{`RANDOM}};
  regs_231_0 = _RAND_231[72:0];
  _RAND_232 = {3{`RANDOM}};
  regs_232_0 = _RAND_232[72:0];
  _RAND_233 = {3{`RANDOM}};
  regs_233_0 = _RAND_233[72:0];
  _RAND_234 = {3{`RANDOM}};
  regs_234_0 = _RAND_234[72:0];
  _RAND_235 = {3{`RANDOM}};
  regs_235_0 = _RAND_235[72:0];
  _RAND_236 = {3{`RANDOM}};
  regs_236_0 = _RAND_236[72:0];
  _RAND_237 = {3{`RANDOM}};
  regs_237_0 = _RAND_237[72:0];
  _RAND_238 = {3{`RANDOM}};
  regs_238_0 = _RAND_238[72:0];
  _RAND_239 = {3{`RANDOM}};
  regs_239_0 = _RAND_239[72:0];
  _RAND_240 = {3{`RANDOM}};
  regs_240_0 = _RAND_240[72:0];
  _RAND_241 = {3{`RANDOM}};
  regs_241_0 = _RAND_241[72:0];
  _RAND_242 = {3{`RANDOM}};
  regs_242_0 = _RAND_242[72:0];
  _RAND_243 = {3{`RANDOM}};
  regs_243_0 = _RAND_243[72:0];
  _RAND_244 = {3{`RANDOM}};
  regs_244_0 = _RAND_244[72:0];
  _RAND_245 = {3{`RANDOM}};
  regs_245_0 = _RAND_245[72:0];
  _RAND_246 = {3{`RANDOM}};
  regs_246_0 = _RAND_246[72:0];
  _RAND_247 = {3{`RANDOM}};
  regs_247_0 = _RAND_247[72:0];
  _RAND_248 = {3{`RANDOM}};
  regs_248_0 = _RAND_248[72:0];
  _RAND_249 = {3{`RANDOM}};
  regs_249_0 = _RAND_249[72:0];
  _RAND_250 = {3{`RANDOM}};
  regs_250_0 = _RAND_250[72:0];
  _RAND_251 = {3{`RANDOM}};
  regs_251_0 = _RAND_251[72:0];
  _RAND_252 = {3{`RANDOM}};
  regs_252_0 = _RAND_252[72:0];
  _RAND_253 = {3{`RANDOM}};
  regs_253_0 = _RAND_253[72:0];
  _RAND_254 = {3{`RANDOM}};
  regs_254_0 = _RAND_254[72:0];
  _RAND_255 = {3{`RANDOM}};
  regs_255_0 = _RAND_255[72:0];
  _RAND_256 = {3{`RANDOM}};
  regs_256_0 = _RAND_256[72:0];
  _RAND_257 = {3{`RANDOM}};
  regs_257_0 = _RAND_257[72:0];
  _RAND_258 = {3{`RANDOM}};
  regs_258_0 = _RAND_258[72:0];
  _RAND_259 = {3{`RANDOM}};
  regs_259_0 = _RAND_259[72:0];
  _RAND_260 = {3{`RANDOM}};
  regs_260_0 = _RAND_260[72:0];
  _RAND_261 = {3{`RANDOM}};
  regs_261_0 = _RAND_261[72:0];
  _RAND_262 = {3{`RANDOM}};
  regs_262_0 = _RAND_262[72:0];
  _RAND_263 = {3{`RANDOM}};
  regs_263_0 = _RAND_263[72:0];
  _RAND_264 = {3{`RANDOM}};
  regs_264_0 = _RAND_264[72:0];
  _RAND_265 = {3{`RANDOM}};
  regs_265_0 = _RAND_265[72:0];
  _RAND_266 = {3{`RANDOM}};
  regs_266_0 = _RAND_266[72:0];
  _RAND_267 = {3{`RANDOM}};
  regs_267_0 = _RAND_267[72:0];
  _RAND_268 = {3{`RANDOM}};
  regs_268_0 = _RAND_268[72:0];
  _RAND_269 = {3{`RANDOM}};
  regs_269_0 = _RAND_269[72:0];
  _RAND_270 = {3{`RANDOM}};
  regs_270_0 = _RAND_270[72:0];
  _RAND_271 = {3{`RANDOM}};
  regs_271_0 = _RAND_271[72:0];
  _RAND_272 = {3{`RANDOM}};
  regs_272_0 = _RAND_272[72:0];
  _RAND_273 = {3{`RANDOM}};
  regs_273_0 = _RAND_273[72:0];
  _RAND_274 = {3{`RANDOM}};
  regs_274_0 = _RAND_274[72:0];
  _RAND_275 = {3{`RANDOM}};
  regs_275_0 = _RAND_275[72:0];
  _RAND_276 = {3{`RANDOM}};
  regs_276_0 = _RAND_276[72:0];
  _RAND_277 = {3{`RANDOM}};
  regs_277_0 = _RAND_277[72:0];
  _RAND_278 = {3{`RANDOM}};
  regs_278_0 = _RAND_278[72:0];
  _RAND_279 = {3{`RANDOM}};
  regs_279_0 = _RAND_279[72:0];
  _RAND_280 = {3{`RANDOM}};
  regs_280_0 = _RAND_280[72:0];
  _RAND_281 = {3{`RANDOM}};
  regs_281_0 = _RAND_281[72:0];
  _RAND_282 = {3{`RANDOM}};
  regs_282_0 = _RAND_282[72:0];
  _RAND_283 = {3{`RANDOM}};
  regs_283_0 = _RAND_283[72:0];
  _RAND_284 = {3{`RANDOM}};
  regs_284_0 = _RAND_284[72:0];
  _RAND_285 = {3{`RANDOM}};
  regs_285_0 = _RAND_285[72:0];
  _RAND_286 = {3{`RANDOM}};
  regs_286_0 = _RAND_286[72:0];
  _RAND_287 = {3{`RANDOM}};
  regs_287_0 = _RAND_287[72:0];
  _RAND_288 = {3{`RANDOM}};
  regs_288_0 = _RAND_288[72:0];
  _RAND_289 = {3{`RANDOM}};
  regs_289_0 = _RAND_289[72:0];
  _RAND_290 = {3{`RANDOM}};
  regs_290_0 = _RAND_290[72:0];
  _RAND_291 = {3{`RANDOM}};
  regs_291_0 = _RAND_291[72:0];
  _RAND_292 = {3{`RANDOM}};
  regs_292_0 = _RAND_292[72:0];
  _RAND_293 = {3{`RANDOM}};
  regs_293_0 = _RAND_293[72:0];
  _RAND_294 = {3{`RANDOM}};
  regs_294_0 = _RAND_294[72:0];
  _RAND_295 = {3{`RANDOM}};
  regs_295_0 = _RAND_295[72:0];
  _RAND_296 = {3{`RANDOM}};
  regs_296_0 = _RAND_296[72:0];
  _RAND_297 = {3{`RANDOM}};
  regs_297_0 = _RAND_297[72:0];
  _RAND_298 = {3{`RANDOM}};
  regs_298_0 = _RAND_298[72:0];
  _RAND_299 = {3{`RANDOM}};
  regs_299_0 = _RAND_299[72:0];
  _RAND_300 = {3{`RANDOM}};
  regs_300_0 = _RAND_300[72:0];
  _RAND_301 = {3{`RANDOM}};
  regs_301_0 = _RAND_301[72:0];
  _RAND_302 = {3{`RANDOM}};
  regs_302_0 = _RAND_302[72:0];
  _RAND_303 = {3{`RANDOM}};
  regs_303_0 = _RAND_303[72:0];
  _RAND_304 = {3{`RANDOM}};
  regs_304_0 = _RAND_304[72:0];
  _RAND_305 = {3{`RANDOM}};
  regs_305_0 = _RAND_305[72:0];
  _RAND_306 = {3{`RANDOM}};
  regs_306_0 = _RAND_306[72:0];
  _RAND_307 = {3{`RANDOM}};
  regs_307_0 = _RAND_307[72:0];
  _RAND_308 = {3{`RANDOM}};
  regs_308_0 = _RAND_308[72:0];
  _RAND_309 = {3{`RANDOM}};
  regs_309_0 = _RAND_309[72:0];
  _RAND_310 = {3{`RANDOM}};
  regs_310_0 = _RAND_310[72:0];
  _RAND_311 = {3{`RANDOM}};
  regs_311_0 = _RAND_311[72:0];
  _RAND_312 = {3{`RANDOM}};
  regs_312_0 = _RAND_312[72:0];
  _RAND_313 = {3{`RANDOM}};
  regs_313_0 = _RAND_313[72:0];
  _RAND_314 = {3{`RANDOM}};
  regs_314_0 = _RAND_314[72:0];
  _RAND_315 = {3{`RANDOM}};
  regs_315_0 = _RAND_315[72:0];
  _RAND_316 = {3{`RANDOM}};
  regs_316_0 = _RAND_316[72:0];
  _RAND_317 = {3{`RANDOM}};
  regs_317_0 = _RAND_317[72:0];
  _RAND_318 = {3{`RANDOM}};
  regs_318_0 = _RAND_318[72:0];
  _RAND_319 = {3{`RANDOM}};
  regs_319_0 = _RAND_319[72:0];
  _RAND_320 = {3{`RANDOM}};
  regs_320_0 = _RAND_320[72:0];
  _RAND_321 = {3{`RANDOM}};
  regs_321_0 = _RAND_321[72:0];
  _RAND_322 = {3{`RANDOM}};
  regs_322_0 = _RAND_322[72:0];
  _RAND_323 = {3{`RANDOM}};
  regs_323_0 = _RAND_323[72:0];
  _RAND_324 = {3{`RANDOM}};
  regs_324_0 = _RAND_324[72:0];
  _RAND_325 = {3{`RANDOM}};
  regs_325_0 = _RAND_325[72:0];
  _RAND_326 = {3{`RANDOM}};
  regs_326_0 = _RAND_326[72:0];
  _RAND_327 = {3{`RANDOM}};
  regs_327_0 = _RAND_327[72:0];
  _RAND_328 = {3{`RANDOM}};
  regs_328_0 = _RAND_328[72:0];
  _RAND_329 = {3{`RANDOM}};
  regs_329_0 = _RAND_329[72:0];
  _RAND_330 = {3{`RANDOM}};
  regs_330_0 = _RAND_330[72:0];
  _RAND_331 = {3{`RANDOM}};
  regs_331_0 = _RAND_331[72:0];
  _RAND_332 = {3{`RANDOM}};
  regs_332_0 = _RAND_332[72:0];
  _RAND_333 = {3{`RANDOM}};
  regs_333_0 = _RAND_333[72:0];
  _RAND_334 = {3{`RANDOM}};
  regs_334_0 = _RAND_334[72:0];
  _RAND_335 = {3{`RANDOM}};
  regs_335_0 = _RAND_335[72:0];
  _RAND_336 = {3{`RANDOM}};
  regs_336_0 = _RAND_336[72:0];
  _RAND_337 = {3{`RANDOM}};
  regs_337_0 = _RAND_337[72:0];
  _RAND_338 = {3{`RANDOM}};
  regs_338_0 = _RAND_338[72:0];
  _RAND_339 = {3{`RANDOM}};
  regs_339_0 = _RAND_339[72:0];
  _RAND_340 = {3{`RANDOM}};
  regs_340_0 = _RAND_340[72:0];
  _RAND_341 = {3{`RANDOM}};
  regs_341_0 = _RAND_341[72:0];
  _RAND_342 = {3{`RANDOM}};
  regs_342_0 = _RAND_342[72:0];
  _RAND_343 = {3{`RANDOM}};
  regs_343_0 = _RAND_343[72:0];
  _RAND_344 = {3{`RANDOM}};
  regs_344_0 = _RAND_344[72:0];
  _RAND_345 = {3{`RANDOM}};
  regs_345_0 = _RAND_345[72:0];
  _RAND_346 = {3{`RANDOM}};
  regs_346_0 = _RAND_346[72:0];
  _RAND_347 = {3{`RANDOM}};
  regs_347_0 = _RAND_347[72:0];
  _RAND_348 = {3{`RANDOM}};
  regs_348_0 = _RAND_348[72:0];
  _RAND_349 = {3{`RANDOM}};
  regs_349_0 = _RAND_349[72:0];
  _RAND_350 = {3{`RANDOM}};
  regs_350_0 = _RAND_350[72:0];
  _RAND_351 = {3{`RANDOM}};
  regs_351_0 = _RAND_351[72:0];
  _RAND_352 = {3{`RANDOM}};
  regs_352_0 = _RAND_352[72:0];
  _RAND_353 = {3{`RANDOM}};
  regs_353_0 = _RAND_353[72:0];
  _RAND_354 = {3{`RANDOM}};
  regs_354_0 = _RAND_354[72:0];
  _RAND_355 = {3{`RANDOM}};
  regs_355_0 = _RAND_355[72:0];
  _RAND_356 = {3{`RANDOM}};
  regs_356_0 = _RAND_356[72:0];
  _RAND_357 = {3{`RANDOM}};
  regs_357_0 = _RAND_357[72:0];
  _RAND_358 = {3{`RANDOM}};
  regs_358_0 = _RAND_358[72:0];
  _RAND_359 = {3{`RANDOM}};
  regs_359_0 = _RAND_359[72:0];
  _RAND_360 = {3{`RANDOM}};
  regs_360_0 = _RAND_360[72:0];
  _RAND_361 = {3{`RANDOM}};
  regs_361_0 = _RAND_361[72:0];
  _RAND_362 = {3{`RANDOM}};
  regs_362_0 = _RAND_362[72:0];
  _RAND_363 = {3{`RANDOM}};
  regs_363_0 = _RAND_363[72:0];
  _RAND_364 = {3{`RANDOM}};
  regs_364_0 = _RAND_364[72:0];
  _RAND_365 = {3{`RANDOM}};
  regs_365_0 = _RAND_365[72:0];
  _RAND_366 = {3{`RANDOM}};
  regs_366_0 = _RAND_366[72:0];
  _RAND_367 = {3{`RANDOM}};
  regs_367_0 = _RAND_367[72:0];
  _RAND_368 = {3{`RANDOM}};
  regs_368_0 = _RAND_368[72:0];
  _RAND_369 = {3{`RANDOM}};
  regs_369_0 = _RAND_369[72:0];
  _RAND_370 = {3{`RANDOM}};
  regs_370_0 = _RAND_370[72:0];
  _RAND_371 = {3{`RANDOM}};
  regs_371_0 = _RAND_371[72:0];
  _RAND_372 = {3{`RANDOM}};
  regs_372_0 = _RAND_372[72:0];
  _RAND_373 = {3{`RANDOM}};
  regs_373_0 = _RAND_373[72:0];
  _RAND_374 = {3{`RANDOM}};
  regs_374_0 = _RAND_374[72:0];
  _RAND_375 = {3{`RANDOM}};
  regs_375_0 = _RAND_375[72:0];
  _RAND_376 = {3{`RANDOM}};
  regs_376_0 = _RAND_376[72:0];
  _RAND_377 = {3{`RANDOM}};
  regs_377_0 = _RAND_377[72:0];
  _RAND_378 = {3{`RANDOM}};
  regs_378_0 = _RAND_378[72:0];
  _RAND_379 = {3{`RANDOM}};
  regs_379_0 = _RAND_379[72:0];
  _RAND_380 = {3{`RANDOM}};
  regs_380_0 = _RAND_380[72:0];
  _RAND_381 = {3{`RANDOM}};
  regs_381_0 = _RAND_381[72:0];
  _RAND_382 = {3{`RANDOM}};
  regs_382_0 = _RAND_382[72:0];
  _RAND_383 = {3{`RANDOM}};
  regs_383_0 = _RAND_383[72:0];
  _RAND_384 = {3{`RANDOM}};
  regs_384_0 = _RAND_384[72:0];
  _RAND_385 = {3{`RANDOM}};
  regs_385_0 = _RAND_385[72:0];
  _RAND_386 = {3{`RANDOM}};
  regs_386_0 = _RAND_386[72:0];
  _RAND_387 = {3{`RANDOM}};
  regs_387_0 = _RAND_387[72:0];
  _RAND_388 = {3{`RANDOM}};
  regs_388_0 = _RAND_388[72:0];
  _RAND_389 = {3{`RANDOM}};
  regs_389_0 = _RAND_389[72:0];
  _RAND_390 = {3{`RANDOM}};
  regs_390_0 = _RAND_390[72:0];
  _RAND_391 = {3{`RANDOM}};
  regs_391_0 = _RAND_391[72:0];
  _RAND_392 = {3{`RANDOM}};
  regs_392_0 = _RAND_392[72:0];
  _RAND_393 = {3{`RANDOM}};
  regs_393_0 = _RAND_393[72:0];
  _RAND_394 = {3{`RANDOM}};
  regs_394_0 = _RAND_394[72:0];
  _RAND_395 = {3{`RANDOM}};
  regs_395_0 = _RAND_395[72:0];
  _RAND_396 = {3{`RANDOM}};
  regs_396_0 = _RAND_396[72:0];
  _RAND_397 = {3{`RANDOM}};
  regs_397_0 = _RAND_397[72:0];
  _RAND_398 = {3{`RANDOM}};
  regs_398_0 = _RAND_398[72:0];
  _RAND_399 = {3{`RANDOM}};
  regs_399_0 = _RAND_399[72:0];
  _RAND_400 = {3{`RANDOM}};
  regs_400_0 = _RAND_400[72:0];
  _RAND_401 = {3{`RANDOM}};
  regs_401_0 = _RAND_401[72:0];
  _RAND_402 = {3{`RANDOM}};
  regs_402_0 = _RAND_402[72:0];
  _RAND_403 = {3{`RANDOM}};
  regs_403_0 = _RAND_403[72:0];
  _RAND_404 = {3{`RANDOM}};
  regs_404_0 = _RAND_404[72:0];
  _RAND_405 = {3{`RANDOM}};
  regs_405_0 = _RAND_405[72:0];
  _RAND_406 = {3{`RANDOM}};
  regs_406_0 = _RAND_406[72:0];
  _RAND_407 = {3{`RANDOM}};
  regs_407_0 = _RAND_407[72:0];
  _RAND_408 = {3{`RANDOM}};
  regs_408_0 = _RAND_408[72:0];
  _RAND_409 = {3{`RANDOM}};
  regs_409_0 = _RAND_409[72:0];
  _RAND_410 = {3{`RANDOM}};
  regs_410_0 = _RAND_410[72:0];
  _RAND_411 = {3{`RANDOM}};
  regs_411_0 = _RAND_411[72:0];
  _RAND_412 = {3{`RANDOM}};
  regs_412_0 = _RAND_412[72:0];
  _RAND_413 = {3{`RANDOM}};
  regs_413_0 = _RAND_413[72:0];
  _RAND_414 = {3{`RANDOM}};
  regs_414_0 = _RAND_414[72:0];
  _RAND_415 = {3{`RANDOM}};
  regs_415_0 = _RAND_415[72:0];
  _RAND_416 = {3{`RANDOM}};
  regs_416_0 = _RAND_416[72:0];
  _RAND_417 = {3{`RANDOM}};
  regs_417_0 = _RAND_417[72:0];
  _RAND_418 = {3{`RANDOM}};
  regs_418_0 = _RAND_418[72:0];
  _RAND_419 = {3{`RANDOM}};
  regs_419_0 = _RAND_419[72:0];
  _RAND_420 = {3{`RANDOM}};
  regs_420_0 = _RAND_420[72:0];
  _RAND_421 = {3{`RANDOM}};
  regs_421_0 = _RAND_421[72:0];
  _RAND_422 = {3{`RANDOM}};
  regs_422_0 = _RAND_422[72:0];
  _RAND_423 = {3{`RANDOM}};
  regs_423_0 = _RAND_423[72:0];
  _RAND_424 = {3{`RANDOM}};
  regs_424_0 = _RAND_424[72:0];
  _RAND_425 = {3{`RANDOM}};
  regs_425_0 = _RAND_425[72:0];
  _RAND_426 = {3{`RANDOM}};
  regs_426_0 = _RAND_426[72:0];
  _RAND_427 = {3{`RANDOM}};
  regs_427_0 = _RAND_427[72:0];
  _RAND_428 = {3{`RANDOM}};
  regs_428_0 = _RAND_428[72:0];
  _RAND_429 = {3{`RANDOM}};
  regs_429_0 = _RAND_429[72:0];
  _RAND_430 = {3{`RANDOM}};
  regs_430_0 = _RAND_430[72:0];
  _RAND_431 = {3{`RANDOM}};
  regs_431_0 = _RAND_431[72:0];
  _RAND_432 = {3{`RANDOM}};
  regs_432_0 = _RAND_432[72:0];
  _RAND_433 = {3{`RANDOM}};
  regs_433_0 = _RAND_433[72:0];
  _RAND_434 = {3{`RANDOM}};
  regs_434_0 = _RAND_434[72:0];
  _RAND_435 = {3{`RANDOM}};
  regs_435_0 = _RAND_435[72:0];
  _RAND_436 = {3{`RANDOM}};
  regs_436_0 = _RAND_436[72:0];
  _RAND_437 = {3{`RANDOM}};
  regs_437_0 = _RAND_437[72:0];
  _RAND_438 = {3{`RANDOM}};
  regs_438_0 = _RAND_438[72:0];
  _RAND_439 = {3{`RANDOM}};
  regs_439_0 = _RAND_439[72:0];
  _RAND_440 = {3{`RANDOM}};
  regs_440_0 = _RAND_440[72:0];
  _RAND_441 = {3{`RANDOM}};
  regs_441_0 = _RAND_441[72:0];
  _RAND_442 = {3{`RANDOM}};
  regs_442_0 = _RAND_442[72:0];
  _RAND_443 = {3{`RANDOM}};
  regs_443_0 = _RAND_443[72:0];
  _RAND_444 = {3{`RANDOM}};
  regs_444_0 = _RAND_444[72:0];
  _RAND_445 = {3{`RANDOM}};
  regs_445_0 = _RAND_445[72:0];
  _RAND_446 = {3{`RANDOM}};
  regs_446_0 = _RAND_446[72:0];
  _RAND_447 = {3{`RANDOM}};
  regs_447_0 = _RAND_447[72:0];
  _RAND_448 = {3{`RANDOM}};
  regs_448_0 = _RAND_448[72:0];
  _RAND_449 = {3{`RANDOM}};
  regs_449_0 = _RAND_449[72:0];
  _RAND_450 = {3{`RANDOM}};
  regs_450_0 = _RAND_450[72:0];
  _RAND_451 = {3{`RANDOM}};
  regs_451_0 = _RAND_451[72:0];
  _RAND_452 = {3{`RANDOM}};
  regs_452_0 = _RAND_452[72:0];
  _RAND_453 = {3{`RANDOM}};
  regs_453_0 = _RAND_453[72:0];
  _RAND_454 = {3{`RANDOM}};
  regs_454_0 = _RAND_454[72:0];
  _RAND_455 = {3{`RANDOM}};
  regs_455_0 = _RAND_455[72:0];
  _RAND_456 = {3{`RANDOM}};
  regs_456_0 = _RAND_456[72:0];
  _RAND_457 = {3{`RANDOM}};
  regs_457_0 = _RAND_457[72:0];
  _RAND_458 = {3{`RANDOM}};
  regs_458_0 = _RAND_458[72:0];
  _RAND_459 = {3{`RANDOM}};
  regs_459_0 = _RAND_459[72:0];
  _RAND_460 = {3{`RANDOM}};
  regs_460_0 = _RAND_460[72:0];
  _RAND_461 = {3{`RANDOM}};
  regs_461_0 = _RAND_461[72:0];
  _RAND_462 = {3{`RANDOM}};
  regs_462_0 = _RAND_462[72:0];
  _RAND_463 = {3{`RANDOM}};
  regs_463_0 = _RAND_463[72:0];
  _RAND_464 = {3{`RANDOM}};
  regs_464_0 = _RAND_464[72:0];
  _RAND_465 = {3{`RANDOM}};
  regs_465_0 = _RAND_465[72:0];
  _RAND_466 = {3{`RANDOM}};
  regs_466_0 = _RAND_466[72:0];
  _RAND_467 = {3{`RANDOM}};
  regs_467_0 = _RAND_467[72:0];
  _RAND_468 = {3{`RANDOM}};
  regs_468_0 = _RAND_468[72:0];
  _RAND_469 = {3{`RANDOM}};
  regs_469_0 = _RAND_469[72:0];
  _RAND_470 = {3{`RANDOM}};
  regs_470_0 = _RAND_470[72:0];
  _RAND_471 = {3{`RANDOM}};
  regs_471_0 = _RAND_471[72:0];
  _RAND_472 = {3{`RANDOM}};
  regs_472_0 = _RAND_472[72:0];
  _RAND_473 = {3{`RANDOM}};
  regs_473_0 = _RAND_473[72:0];
  _RAND_474 = {3{`RANDOM}};
  regs_474_0 = _RAND_474[72:0];
  _RAND_475 = {3{`RANDOM}};
  regs_475_0 = _RAND_475[72:0];
  _RAND_476 = {3{`RANDOM}};
  regs_476_0 = _RAND_476[72:0];
  _RAND_477 = {3{`RANDOM}};
  regs_477_0 = _RAND_477[72:0];
  _RAND_478 = {3{`RANDOM}};
  regs_478_0 = _RAND_478[72:0];
  _RAND_479 = {3{`RANDOM}};
  regs_479_0 = _RAND_479[72:0];
  _RAND_480 = {3{`RANDOM}};
  regs_480_0 = _RAND_480[72:0];
  _RAND_481 = {3{`RANDOM}};
  regs_481_0 = _RAND_481[72:0];
  _RAND_482 = {3{`RANDOM}};
  regs_482_0 = _RAND_482[72:0];
  _RAND_483 = {3{`RANDOM}};
  regs_483_0 = _RAND_483[72:0];
  _RAND_484 = {3{`RANDOM}};
  regs_484_0 = _RAND_484[72:0];
  _RAND_485 = {3{`RANDOM}};
  regs_485_0 = _RAND_485[72:0];
  _RAND_486 = {3{`RANDOM}};
  regs_486_0 = _RAND_486[72:0];
  _RAND_487 = {3{`RANDOM}};
  regs_487_0 = _RAND_487[72:0];
  _RAND_488 = {3{`RANDOM}};
  regs_488_0 = _RAND_488[72:0];
  _RAND_489 = {3{`RANDOM}};
  regs_489_0 = _RAND_489[72:0];
  _RAND_490 = {3{`RANDOM}};
  regs_490_0 = _RAND_490[72:0];
  _RAND_491 = {3{`RANDOM}};
  regs_491_0 = _RAND_491[72:0];
  _RAND_492 = {3{`RANDOM}};
  regs_492_0 = _RAND_492[72:0];
  _RAND_493 = {3{`RANDOM}};
  regs_493_0 = _RAND_493[72:0];
  _RAND_494 = {3{`RANDOM}};
  regs_494_0 = _RAND_494[72:0];
  _RAND_495 = {3{`RANDOM}};
  regs_495_0 = _RAND_495[72:0];
  _RAND_496 = {3{`RANDOM}};
  regs_496_0 = _RAND_496[72:0];
  _RAND_497 = {3{`RANDOM}};
  regs_497_0 = _RAND_497[72:0];
  _RAND_498 = {3{`RANDOM}};
  regs_498_0 = _RAND_498[72:0];
  _RAND_499 = {3{`RANDOM}};
  regs_499_0 = _RAND_499[72:0];
  _RAND_500 = {3{`RANDOM}};
  regs_500_0 = _RAND_500[72:0];
  _RAND_501 = {3{`RANDOM}};
  regs_501_0 = _RAND_501[72:0];
  _RAND_502 = {3{`RANDOM}};
  regs_502_0 = _RAND_502[72:0];
  _RAND_503 = {3{`RANDOM}};
  regs_503_0 = _RAND_503[72:0];
  _RAND_504 = {3{`RANDOM}};
  regs_504_0 = _RAND_504[72:0];
  _RAND_505 = {3{`RANDOM}};
  regs_505_0 = _RAND_505[72:0];
  _RAND_506 = {3{`RANDOM}};
  regs_506_0 = _RAND_506[72:0];
  _RAND_507 = {3{`RANDOM}};
  regs_507_0 = _RAND_507[72:0];
  _RAND_508 = {3{`RANDOM}};
  regs_508_0 = _RAND_508[72:0];
  _RAND_509 = {3{`RANDOM}};
  regs_509_0 = _RAND_509[72:0];
  _RAND_510 = {3{`RANDOM}};
  regs_510_0 = _RAND_510[72:0];
  _RAND_511 = {3{`RANDOM}};
  regs_511_0 = _RAND_511[72:0];
  _RAND_512 = {1{`RANDOM}};
  resetState = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  resetSet = _RAND_513[8:0];
  _RAND_514 = {3{`RANDOM}};
  rdata_r_0 = _RAND_514[72:0];
  _RAND_515 = {1{`RANDOM}};
  rdata_REG = _RAND_515[0:0];
  _RAND_516 = {3{`RANDOM}};
  rdata_r_1_0 = _RAND_516[72:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BPU_inorder(
  input         clock,
  input         reset,
  input         io_in_pc_valid, // @[src/main/scala/nutcore/frontend/BPU.scala 281:14]
  input  [38:0] io_in_pc_bits, // @[src/main/scala/nutcore/frontend/BPU.scala 281:14]
  output [38:0] io_out_target, // @[src/main/scala/nutcore/frontend/BPU.scala 281:14]
  output        io_out_valid, // @[src/main/scala/nutcore/frontend/BPU.scala 281:14]
  input         io_flush, // @[src/main/scala/nutcore/frontend/BPU.scala 281:14]
  output [2:0]  io_brIdx, // @[src/main/scala/nutcore/frontend/BPU.scala 281:14]
  output        io_crosslineJump, // @[src/main/scala/nutcore/frontend/BPU.scala 281:14]
  input         MOUFlushICache,
  input         bpuUpdateReq_valid,
  input  [38:0] bpuUpdateReq_pc,
  input         bpuUpdateReq_isMissPredict,
  input  [38:0] bpuUpdateReq_actualTarget,
  input         bpuUpdateReq_actualTaken,
  input  [6:0]  bpuUpdateReq_fuOpType,
  input  [1:0]  bpuUpdateReq_btbType,
  input         bpuUpdateReq_isRVC,
  input         MOUFlushTLB
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [63:0] _RAND_516;
  reg [63:0] _RAND_517;
  reg [63:0] _RAND_518;
  reg [63:0] _RAND_519;
  reg [63:0] _RAND_520;
  reg [63:0] _RAND_521;
  reg [63:0] _RAND_522;
  reg [63:0] _RAND_523;
  reg [63:0] _RAND_524;
  reg [63:0] _RAND_525;
  reg [63:0] _RAND_526;
  reg [63:0] _RAND_527;
  reg [63:0] _RAND_528;
  reg [63:0] _RAND_529;
  reg [63:0] _RAND_530;
  reg [63:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [63:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [63:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
`endif // RANDOMIZE_REG_INIT
  wire  btb_clock; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire  btb_reset; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire  btb_io_r_req_ready; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire  btb_io_r_req_valid; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [8:0] btb_io_r_req_bits_setIdx; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [27:0] btb_io_r_resp_data_0_tag; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [1:0] btb_io_r_resp_data_0__type; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [38:0] btb_io_r_resp_data_0_target; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [2:0] btb_io_r_resp_data_0_brIdx; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire  btb_io_r_resp_data_0_valid; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire  btb_io_w_req_valid; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [8:0] btb_io_w_req_bits_setIdx; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [27:0] btb_io_w_req_bits_data_tag; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [1:0] btb_io_w_req_bits_data__type; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [38:0] btb_io_w_req_bits_data_target; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [2:0] btb_io_w_req_bits_data_brIdx; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  reg  flush; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_0 = io_in_pc_valid ? 1'h0 : flush; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_1 = io_flush | _GEN_0; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg [38:0] pcLatch; // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
  wire [27:0] btbRead_tag = btb_io_r_resp_data_0_tag; // @[src/main/scala/nutcore/frontend/BPU.scala 315:21 316:11]
  wire  btbRead_valid = btb_io_r_resp_data_0_valid; // @[src/main/scala/nutcore/frontend/BPU.scala 315:21 316:11]
  wire  _btbHit_T_7 = btb_io_r_req_ready & btb_io_r_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  btbHit_REG; // @[src/main/scala/nutcore/frontend/BPU.scala 320:93]
  wire [2:0] btbRead_brIdx = btb_io_r_resp_data_0_brIdx; // @[src/main/scala/nutcore/frontend/BPU.scala 315:21 316:11]
  wire  btbHit = btbRead_valid & btbRead_tag == pcLatch[38:11] & ~flush & btbHit_REG & ~(pcLatch[1] & btbRead_brIdx[0]); // @[src/main/scala/nutcore/frontend/BPU.scala 320:129]
  wire  crosslineJump = btbRead_brIdx[2] & btbHit; // @[src/main/scala/nutcore/frontend/BPU.scala 327:40]
  wire [1:0] _T_20 = io_out_valid ? 2'h3 : 2'h0; // @[src/main/scala/nutcore/frontend/BPU.scala 332:94]
  reg [1:0] regs__0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__1; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__2; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__3; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__4; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__5; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__6; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__7; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__8; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__9; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__10; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__11; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__12; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__13; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__14; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__15; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__16; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__17; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__18; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__19; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__20; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__21; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__22; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__23; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__24; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__25; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__26; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__27; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__28; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__29; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__30; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__31; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__32; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__33; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__34; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__35; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__36; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__37; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__38; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__39; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__40; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__41; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__42; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__43; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__44; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__45; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__46; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__47; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__48; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__49; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__50; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__51; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__52; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__53; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__54; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__55; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__56; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__57; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__58; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__59; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__60; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__61; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__62; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__63; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__64; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__65; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__66; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__67; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__68; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__69; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__70; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__71; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__72; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__73; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__74; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__75; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__76; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__77; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__78; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__79; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__80; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__81; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__82; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__83; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__84; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__85; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__86; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__87; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__88; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__89; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__90; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__91; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__92; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__93; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__94; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__95; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__96; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__97; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__98; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__99; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__100; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__101; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__102; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__103; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__104; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__105; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__106; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__107; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__108; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__109; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__110; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__111; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__112; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__113; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__114; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__115; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__116; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__117; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__118; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__119; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__120; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__121; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__122; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__123; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__124; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__125; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__126; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__127; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__128; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__129; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__130; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__131; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__132; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__133; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__134; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__135; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__136; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__137; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__138; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__139; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__140; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__141; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__142; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__143; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__144; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__145; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__146; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__147; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__148; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__149; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__150; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__151; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__152; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__153; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__154; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__155; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__156; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__157; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__158; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__159; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__160; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__161; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__162; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__163; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__164; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__165; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__166; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__167; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__168; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__169; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__170; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__171; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__172; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__173; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__174; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__175; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__176; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__177; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__178; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__179; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__180; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__181; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__182; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__183; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__184; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__185; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__186; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__187; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__188; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__189; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__190; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__191; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__192; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__193; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__194; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__195; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__196; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__197; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__198; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__199; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__200; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__201; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__202; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__203; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__204; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__205; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__206; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__207; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__208; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__209; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__210; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__211; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__212; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__213; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__214; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__215; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__216; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__217; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__218; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__219; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__220; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__221; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__222; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__223; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__224; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__225; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__226; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__227; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__228; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__229; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__230; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__231; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__232; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__233; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__234; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__235; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__236; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__237; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__238; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__239; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__240; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__241; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__242; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__243; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__244; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__245; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__246; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__247; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__248; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__249; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__250; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__251; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__252; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__253; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__254; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__255; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__256; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__257; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__258; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__259; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__260; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__261; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__262; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__263; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__264; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__265; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__266; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__267; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__268; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__269; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__270; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__271; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__272; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__273; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__274; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__275; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__276; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__277; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__278; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__279; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__280; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__281; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__282; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__283; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__284; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__285; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__286; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__287; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__288; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__289; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__290; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__291; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__292; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__293; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__294; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__295; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__296; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__297; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__298; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__299; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__300; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__301; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__302; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__303; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__304; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__305; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__306; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__307; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__308; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__309; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__310; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__311; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__312; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__313; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__314; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__315; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__316; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__317; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__318; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__319; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__320; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__321; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__322; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__323; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__324; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__325; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__326; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__327; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__328; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__329; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__330; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__331; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__332; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__333; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__334; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__335; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__336; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__337; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__338; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__339; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__340; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__341; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__342; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__343; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__344; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__345; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__346; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__347; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__348; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__349; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__350; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__351; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__352; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__353; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__354; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__355; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__356; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__357; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__358; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__359; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__360; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__361; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__362; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__363; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__364; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__365; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__366; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__367; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__368; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__369; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__370; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__371; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__372; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__373; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__374; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__375; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__376; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__377; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__378; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__379; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__380; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__381; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__382; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__383; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__384; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__385; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__386; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__387; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__388; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__389; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__390; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__391; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__392; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__393; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__394; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__395; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__396; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__397; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__398; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__399; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__400; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__401; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__402; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__403; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__404; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__405; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__406; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__407; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__408; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__409; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__410; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__411; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__412; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__413; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__414; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__415; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__416; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__417; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__418; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__419; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__420; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__421; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__422; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__423; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__424; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__425; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__426; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__427; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__428; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__429; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__430; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__431; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__432; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__433; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__434; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__435; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__436; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__437; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__438; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__439; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__440; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__441; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__442; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__443; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__444; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__445; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__446; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__447; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__448; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__449; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__450; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__451; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__452; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__453; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__454; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__455; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__456; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__457; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__458; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__459; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__460; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__461; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__462; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__463; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__464; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__465; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__466; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__467; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__468; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__469; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__470; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__471; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__472; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__473; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__474; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__475; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__476; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__477; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__478; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__479; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__480; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__481; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__482; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__483; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__484; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__485; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__486; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__487; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__488; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__489; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__490; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__491; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__492; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__493; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__494; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__495; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__496; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__497; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__498; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__499; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__500; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__501; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__502; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__503; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__504; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__505; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__506; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__507; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__508; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__509; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__510; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] regs__511; // @[src/main/scala/utils/RegMem.scala 7:21]
  wire [1:0] _GEN_4 = 9'h1 == io_in_pc_bits[10:2] ? regs__1 : regs__0; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_5 = 9'h2 == io_in_pc_bits[10:2] ? regs__2 : _GEN_4; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_6 = 9'h3 == io_in_pc_bits[10:2] ? regs__3 : _GEN_5; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_7 = 9'h4 == io_in_pc_bits[10:2] ? regs__4 : _GEN_6; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_8 = 9'h5 == io_in_pc_bits[10:2] ? regs__5 : _GEN_7; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_9 = 9'h6 == io_in_pc_bits[10:2] ? regs__6 : _GEN_8; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_10 = 9'h7 == io_in_pc_bits[10:2] ? regs__7 : _GEN_9; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_11 = 9'h8 == io_in_pc_bits[10:2] ? regs__8 : _GEN_10; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_12 = 9'h9 == io_in_pc_bits[10:2] ? regs__9 : _GEN_11; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_13 = 9'ha == io_in_pc_bits[10:2] ? regs__10 : _GEN_12; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_14 = 9'hb == io_in_pc_bits[10:2] ? regs__11 : _GEN_13; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_15 = 9'hc == io_in_pc_bits[10:2] ? regs__12 : _GEN_14; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_16 = 9'hd == io_in_pc_bits[10:2] ? regs__13 : _GEN_15; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_17 = 9'he == io_in_pc_bits[10:2] ? regs__14 : _GEN_16; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_18 = 9'hf == io_in_pc_bits[10:2] ? regs__15 : _GEN_17; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_19 = 9'h10 == io_in_pc_bits[10:2] ? regs__16 : _GEN_18; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_20 = 9'h11 == io_in_pc_bits[10:2] ? regs__17 : _GEN_19; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_21 = 9'h12 == io_in_pc_bits[10:2] ? regs__18 : _GEN_20; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_22 = 9'h13 == io_in_pc_bits[10:2] ? regs__19 : _GEN_21; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_23 = 9'h14 == io_in_pc_bits[10:2] ? regs__20 : _GEN_22; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_24 = 9'h15 == io_in_pc_bits[10:2] ? regs__21 : _GEN_23; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_25 = 9'h16 == io_in_pc_bits[10:2] ? regs__22 : _GEN_24; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_26 = 9'h17 == io_in_pc_bits[10:2] ? regs__23 : _GEN_25; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_27 = 9'h18 == io_in_pc_bits[10:2] ? regs__24 : _GEN_26; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_28 = 9'h19 == io_in_pc_bits[10:2] ? regs__25 : _GEN_27; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_29 = 9'h1a == io_in_pc_bits[10:2] ? regs__26 : _GEN_28; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_30 = 9'h1b == io_in_pc_bits[10:2] ? regs__27 : _GEN_29; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_31 = 9'h1c == io_in_pc_bits[10:2] ? regs__28 : _GEN_30; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_32 = 9'h1d == io_in_pc_bits[10:2] ? regs__29 : _GEN_31; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_33 = 9'h1e == io_in_pc_bits[10:2] ? regs__30 : _GEN_32; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_34 = 9'h1f == io_in_pc_bits[10:2] ? regs__31 : _GEN_33; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_35 = 9'h20 == io_in_pc_bits[10:2] ? regs__32 : _GEN_34; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_36 = 9'h21 == io_in_pc_bits[10:2] ? regs__33 : _GEN_35; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_37 = 9'h22 == io_in_pc_bits[10:2] ? regs__34 : _GEN_36; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_38 = 9'h23 == io_in_pc_bits[10:2] ? regs__35 : _GEN_37; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_39 = 9'h24 == io_in_pc_bits[10:2] ? regs__36 : _GEN_38; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_40 = 9'h25 == io_in_pc_bits[10:2] ? regs__37 : _GEN_39; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_41 = 9'h26 == io_in_pc_bits[10:2] ? regs__38 : _GEN_40; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_42 = 9'h27 == io_in_pc_bits[10:2] ? regs__39 : _GEN_41; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_43 = 9'h28 == io_in_pc_bits[10:2] ? regs__40 : _GEN_42; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_44 = 9'h29 == io_in_pc_bits[10:2] ? regs__41 : _GEN_43; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_45 = 9'h2a == io_in_pc_bits[10:2] ? regs__42 : _GEN_44; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_46 = 9'h2b == io_in_pc_bits[10:2] ? regs__43 : _GEN_45; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_47 = 9'h2c == io_in_pc_bits[10:2] ? regs__44 : _GEN_46; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_48 = 9'h2d == io_in_pc_bits[10:2] ? regs__45 : _GEN_47; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_49 = 9'h2e == io_in_pc_bits[10:2] ? regs__46 : _GEN_48; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_50 = 9'h2f == io_in_pc_bits[10:2] ? regs__47 : _GEN_49; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_51 = 9'h30 == io_in_pc_bits[10:2] ? regs__48 : _GEN_50; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_52 = 9'h31 == io_in_pc_bits[10:2] ? regs__49 : _GEN_51; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_53 = 9'h32 == io_in_pc_bits[10:2] ? regs__50 : _GEN_52; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_54 = 9'h33 == io_in_pc_bits[10:2] ? regs__51 : _GEN_53; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_55 = 9'h34 == io_in_pc_bits[10:2] ? regs__52 : _GEN_54; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_56 = 9'h35 == io_in_pc_bits[10:2] ? regs__53 : _GEN_55; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_57 = 9'h36 == io_in_pc_bits[10:2] ? regs__54 : _GEN_56; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_58 = 9'h37 == io_in_pc_bits[10:2] ? regs__55 : _GEN_57; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_59 = 9'h38 == io_in_pc_bits[10:2] ? regs__56 : _GEN_58; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_60 = 9'h39 == io_in_pc_bits[10:2] ? regs__57 : _GEN_59; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_61 = 9'h3a == io_in_pc_bits[10:2] ? regs__58 : _GEN_60; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_62 = 9'h3b == io_in_pc_bits[10:2] ? regs__59 : _GEN_61; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_63 = 9'h3c == io_in_pc_bits[10:2] ? regs__60 : _GEN_62; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_64 = 9'h3d == io_in_pc_bits[10:2] ? regs__61 : _GEN_63; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_65 = 9'h3e == io_in_pc_bits[10:2] ? regs__62 : _GEN_64; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_66 = 9'h3f == io_in_pc_bits[10:2] ? regs__63 : _GEN_65; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_67 = 9'h40 == io_in_pc_bits[10:2] ? regs__64 : _GEN_66; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_68 = 9'h41 == io_in_pc_bits[10:2] ? regs__65 : _GEN_67; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_69 = 9'h42 == io_in_pc_bits[10:2] ? regs__66 : _GEN_68; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_70 = 9'h43 == io_in_pc_bits[10:2] ? regs__67 : _GEN_69; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_71 = 9'h44 == io_in_pc_bits[10:2] ? regs__68 : _GEN_70; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_72 = 9'h45 == io_in_pc_bits[10:2] ? regs__69 : _GEN_71; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_73 = 9'h46 == io_in_pc_bits[10:2] ? regs__70 : _GEN_72; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_74 = 9'h47 == io_in_pc_bits[10:2] ? regs__71 : _GEN_73; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_75 = 9'h48 == io_in_pc_bits[10:2] ? regs__72 : _GEN_74; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_76 = 9'h49 == io_in_pc_bits[10:2] ? regs__73 : _GEN_75; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_77 = 9'h4a == io_in_pc_bits[10:2] ? regs__74 : _GEN_76; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_78 = 9'h4b == io_in_pc_bits[10:2] ? regs__75 : _GEN_77; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_79 = 9'h4c == io_in_pc_bits[10:2] ? regs__76 : _GEN_78; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_80 = 9'h4d == io_in_pc_bits[10:2] ? regs__77 : _GEN_79; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_81 = 9'h4e == io_in_pc_bits[10:2] ? regs__78 : _GEN_80; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_82 = 9'h4f == io_in_pc_bits[10:2] ? regs__79 : _GEN_81; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_83 = 9'h50 == io_in_pc_bits[10:2] ? regs__80 : _GEN_82; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_84 = 9'h51 == io_in_pc_bits[10:2] ? regs__81 : _GEN_83; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_85 = 9'h52 == io_in_pc_bits[10:2] ? regs__82 : _GEN_84; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_86 = 9'h53 == io_in_pc_bits[10:2] ? regs__83 : _GEN_85; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_87 = 9'h54 == io_in_pc_bits[10:2] ? regs__84 : _GEN_86; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_88 = 9'h55 == io_in_pc_bits[10:2] ? regs__85 : _GEN_87; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_89 = 9'h56 == io_in_pc_bits[10:2] ? regs__86 : _GEN_88; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_90 = 9'h57 == io_in_pc_bits[10:2] ? regs__87 : _GEN_89; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_91 = 9'h58 == io_in_pc_bits[10:2] ? regs__88 : _GEN_90; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_92 = 9'h59 == io_in_pc_bits[10:2] ? regs__89 : _GEN_91; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_93 = 9'h5a == io_in_pc_bits[10:2] ? regs__90 : _GEN_92; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_94 = 9'h5b == io_in_pc_bits[10:2] ? regs__91 : _GEN_93; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_95 = 9'h5c == io_in_pc_bits[10:2] ? regs__92 : _GEN_94; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_96 = 9'h5d == io_in_pc_bits[10:2] ? regs__93 : _GEN_95; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_97 = 9'h5e == io_in_pc_bits[10:2] ? regs__94 : _GEN_96; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_98 = 9'h5f == io_in_pc_bits[10:2] ? regs__95 : _GEN_97; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_99 = 9'h60 == io_in_pc_bits[10:2] ? regs__96 : _GEN_98; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_100 = 9'h61 == io_in_pc_bits[10:2] ? regs__97 : _GEN_99; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_101 = 9'h62 == io_in_pc_bits[10:2] ? regs__98 : _GEN_100; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_102 = 9'h63 == io_in_pc_bits[10:2] ? regs__99 : _GEN_101; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_103 = 9'h64 == io_in_pc_bits[10:2] ? regs__100 : _GEN_102; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_104 = 9'h65 == io_in_pc_bits[10:2] ? regs__101 : _GEN_103; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_105 = 9'h66 == io_in_pc_bits[10:2] ? regs__102 : _GEN_104; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_106 = 9'h67 == io_in_pc_bits[10:2] ? regs__103 : _GEN_105; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_107 = 9'h68 == io_in_pc_bits[10:2] ? regs__104 : _GEN_106; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_108 = 9'h69 == io_in_pc_bits[10:2] ? regs__105 : _GEN_107; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_109 = 9'h6a == io_in_pc_bits[10:2] ? regs__106 : _GEN_108; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_110 = 9'h6b == io_in_pc_bits[10:2] ? regs__107 : _GEN_109; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_111 = 9'h6c == io_in_pc_bits[10:2] ? regs__108 : _GEN_110; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_112 = 9'h6d == io_in_pc_bits[10:2] ? regs__109 : _GEN_111; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_113 = 9'h6e == io_in_pc_bits[10:2] ? regs__110 : _GEN_112; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_114 = 9'h6f == io_in_pc_bits[10:2] ? regs__111 : _GEN_113; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_115 = 9'h70 == io_in_pc_bits[10:2] ? regs__112 : _GEN_114; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_116 = 9'h71 == io_in_pc_bits[10:2] ? regs__113 : _GEN_115; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_117 = 9'h72 == io_in_pc_bits[10:2] ? regs__114 : _GEN_116; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_118 = 9'h73 == io_in_pc_bits[10:2] ? regs__115 : _GEN_117; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_119 = 9'h74 == io_in_pc_bits[10:2] ? regs__116 : _GEN_118; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_120 = 9'h75 == io_in_pc_bits[10:2] ? regs__117 : _GEN_119; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_121 = 9'h76 == io_in_pc_bits[10:2] ? regs__118 : _GEN_120; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_122 = 9'h77 == io_in_pc_bits[10:2] ? regs__119 : _GEN_121; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_123 = 9'h78 == io_in_pc_bits[10:2] ? regs__120 : _GEN_122; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_124 = 9'h79 == io_in_pc_bits[10:2] ? regs__121 : _GEN_123; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_125 = 9'h7a == io_in_pc_bits[10:2] ? regs__122 : _GEN_124; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_126 = 9'h7b == io_in_pc_bits[10:2] ? regs__123 : _GEN_125; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_127 = 9'h7c == io_in_pc_bits[10:2] ? regs__124 : _GEN_126; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_128 = 9'h7d == io_in_pc_bits[10:2] ? regs__125 : _GEN_127; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_129 = 9'h7e == io_in_pc_bits[10:2] ? regs__126 : _GEN_128; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_130 = 9'h7f == io_in_pc_bits[10:2] ? regs__127 : _GEN_129; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_131 = 9'h80 == io_in_pc_bits[10:2] ? regs__128 : _GEN_130; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_132 = 9'h81 == io_in_pc_bits[10:2] ? regs__129 : _GEN_131; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_133 = 9'h82 == io_in_pc_bits[10:2] ? regs__130 : _GEN_132; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_134 = 9'h83 == io_in_pc_bits[10:2] ? regs__131 : _GEN_133; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_135 = 9'h84 == io_in_pc_bits[10:2] ? regs__132 : _GEN_134; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_136 = 9'h85 == io_in_pc_bits[10:2] ? regs__133 : _GEN_135; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_137 = 9'h86 == io_in_pc_bits[10:2] ? regs__134 : _GEN_136; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_138 = 9'h87 == io_in_pc_bits[10:2] ? regs__135 : _GEN_137; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_139 = 9'h88 == io_in_pc_bits[10:2] ? regs__136 : _GEN_138; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_140 = 9'h89 == io_in_pc_bits[10:2] ? regs__137 : _GEN_139; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_141 = 9'h8a == io_in_pc_bits[10:2] ? regs__138 : _GEN_140; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_142 = 9'h8b == io_in_pc_bits[10:2] ? regs__139 : _GEN_141; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_143 = 9'h8c == io_in_pc_bits[10:2] ? regs__140 : _GEN_142; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_144 = 9'h8d == io_in_pc_bits[10:2] ? regs__141 : _GEN_143; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_145 = 9'h8e == io_in_pc_bits[10:2] ? regs__142 : _GEN_144; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_146 = 9'h8f == io_in_pc_bits[10:2] ? regs__143 : _GEN_145; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_147 = 9'h90 == io_in_pc_bits[10:2] ? regs__144 : _GEN_146; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_148 = 9'h91 == io_in_pc_bits[10:2] ? regs__145 : _GEN_147; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_149 = 9'h92 == io_in_pc_bits[10:2] ? regs__146 : _GEN_148; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_150 = 9'h93 == io_in_pc_bits[10:2] ? regs__147 : _GEN_149; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_151 = 9'h94 == io_in_pc_bits[10:2] ? regs__148 : _GEN_150; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_152 = 9'h95 == io_in_pc_bits[10:2] ? regs__149 : _GEN_151; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_153 = 9'h96 == io_in_pc_bits[10:2] ? regs__150 : _GEN_152; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_154 = 9'h97 == io_in_pc_bits[10:2] ? regs__151 : _GEN_153; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_155 = 9'h98 == io_in_pc_bits[10:2] ? regs__152 : _GEN_154; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_156 = 9'h99 == io_in_pc_bits[10:2] ? regs__153 : _GEN_155; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_157 = 9'h9a == io_in_pc_bits[10:2] ? regs__154 : _GEN_156; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_158 = 9'h9b == io_in_pc_bits[10:2] ? regs__155 : _GEN_157; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_159 = 9'h9c == io_in_pc_bits[10:2] ? regs__156 : _GEN_158; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_160 = 9'h9d == io_in_pc_bits[10:2] ? regs__157 : _GEN_159; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_161 = 9'h9e == io_in_pc_bits[10:2] ? regs__158 : _GEN_160; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_162 = 9'h9f == io_in_pc_bits[10:2] ? regs__159 : _GEN_161; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_163 = 9'ha0 == io_in_pc_bits[10:2] ? regs__160 : _GEN_162; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_164 = 9'ha1 == io_in_pc_bits[10:2] ? regs__161 : _GEN_163; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_165 = 9'ha2 == io_in_pc_bits[10:2] ? regs__162 : _GEN_164; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_166 = 9'ha3 == io_in_pc_bits[10:2] ? regs__163 : _GEN_165; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_167 = 9'ha4 == io_in_pc_bits[10:2] ? regs__164 : _GEN_166; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_168 = 9'ha5 == io_in_pc_bits[10:2] ? regs__165 : _GEN_167; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_169 = 9'ha6 == io_in_pc_bits[10:2] ? regs__166 : _GEN_168; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_170 = 9'ha7 == io_in_pc_bits[10:2] ? regs__167 : _GEN_169; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_171 = 9'ha8 == io_in_pc_bits[10:2] ? regs__168 : _GEN_170; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_172 = 9'ha9 == io_in_pc_bits[10:2] ? regs__169 : _GEN_171; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_173 = 9'haa == io_in_pc_bits[10:2] ? regs__170 : _GEN_172; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_174 = 9'hab == io_in_pc_bits[10:2] ? regs__171 : _GEN_173; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_175 = 9'hac == io_in_pc_bits[10:2] ? regs__172 : _GEN_174; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_176 = 9'had == io_in_pc_bits[10:2] ? regs__173 : _GEN_175; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_177 = 9'hae == io_in_pc_bits[10:2] ? regs__174 : _GEN_176; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_178 = 9'haf == io_in_pc_bits[10:2] ? regs__175 : _GEN_177; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_179 = 9'hb0 == io_in_pc_bits[10:2] ? regs__176 : _GEN_178; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_180 = 9'hb1 == io_in_pc_bits[10:2] ? regs__177 : _GEN_179; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_181 = 9'hb2 == io_in_pc_bits[10:2] ? regs__178 : _GEN_180; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_182 = 9'hb3 == io_in_pc_bits[10:2] ? regs__179 : _GEN_181; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_183 = 9'hb4 == io_in_pc_bits[10:2] ? regs__180 : _GEN_182; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_184 = 9'hb5 == io_in_pc_bits[10:2] ? regs__181 : _GEN_183; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_185 = 9'hb6 == io_in_pc_bits[10:2] ? regs__182 : _GEN_184; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_186 = 9'hb7 == io_in_pc_bits[10:2] ? regs__183 : _GEN_185; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_187 = 9'hb8 == io_in_pc_bits[10:2] ? regs__184 : _GEN_186; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_188 = 9'hb9 == io_in_pc_bits[10:2] ? regs__185 : _GEN_187; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_189 = 9'hba == io_in_pc_bits[10:2] ? regs__186 : _GEN_188; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_190 = 9'hbb == io_in_pc_bits[10:2] ? regs__187 : _GEN_189; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_191 = 9'hbc == io_in_pc_bits[10:2] ? regs__188 : _GEN_190; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_192 = 9'hbd == io_in_pc_bits[10:2] ? regs__189 : _GEN_191; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_193 = 9'hbe == io_in_pc_bits[10:2] ? regs__190 : _GEN_192; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_194 = 9'hbf == io_in_pc_bits[10:2] ? regs__191 : _GEN_193; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_195 = 9'hc0 == io_in_pc_bits[10:2] ? regs__192 : _GEN_194; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_196 = 9'hc1 == io_in_pc_bits[10:2] ? regs__193 : _GEN_195; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_197 = 9'hc2 == io_in_pc_bits[10:2] ? regs__194 : _GEN_196; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_198 = 9'hc3 == io_in_pc_bits[10:2] ? regs__195 : _GEN_197; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_199 = 9'hc4 == io_in_pc_bits[10:2] ? regs__196 : _GEN_198; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_200 = 9'hc5 == io_in_pc_bits[10:2] ? regs__197 : _GEN_199; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_201 = 9'hc6 == io_in_pc_bits[10:2] ? regs__198 : _GEN_200; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_202 = 9'hc7 == io_in_pc_bits[10:2] ? regs__199 : _GEN_201; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_203 = 9'hc8 == io_in_pc_bits[10:2] ? regs__200 : _GEN_202; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_204 = 9'hc9 == io_in_pc_bits[10:2] ? regs__201 : _GEN_203; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_205 = 9'hca == io_in_pc_bits[10:2] ? regs__202 : _GEN_204; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_206 = 9'hcb == io_in_pc_bits[10:2] ? regs__203 : _GEN_205; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_207 = 9'hcc == io_in_pc_bits[10:2] ? regs__204 : _GEN_206; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_208 = 9'hcd == io_in_pc_bits[10:2] ? regs__205 : _GEN_207; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_209 = 9'hce == io_in_pc_bits[10:2] ? regs__206 : _GEN_208; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_210 = 9'hcf == io_in_pc_bits[10:2] ? regs__207 : _GEN_209; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_211 = 9'hd0 == io_in_pc_bits[10:2] ? regs__208 : _GEN_210; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_212 = 9'hd1 == io_in_pc_bits[10:2] ? regs__209 : _GEN_211; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_213 = 9'hd2 == io_in_pc_bits[10:2] ? regs__210 : _GEN_212; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_214 = 9'hd3 == io_in_pc_bits[10:2] ? regs__211 : _GEN_213; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_215 = 9'hd4 == io_in_pc_bits[10:2] ? regs__212 : _GEN_214; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_216 = 9'hd5 == io_in_pc_bits[10:2] ? regs__213 : _GEN_215; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_217 = 9'hd6 == io_in_pc_bits[10:2] ? regs__214 : _GEN_216; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_218 = 9'hd7 == io_in_pc_bits[10:2] ? regs__215 : _GEN_217; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_219 = 9'hd8 == io_in_pc_bits[10:2] ? regs__216 : _GEN_218; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_220 = 9'hd9 == io_in_pc_bits[10:2] ? regs__217 : _GEN_219; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_221 = 9'hda == io_in_pc_bits[10:2] ? regs__218 : _GEN_220; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_222 = 9'hdb == io_in_pc_bits[10:2] ? regs__219 : _GEN_221; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_223 = 9'hdc == io_in_pc_bits[10:2] ? regs__220 : _GEN_222; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_224 = 9'hdd == io_in_pc_bits[10:2] ? regs__221 : _GEN_223; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_225 = 9'hde == io_in_pc_bits[10:2] ? regs__222 : _GEN_224; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_226 = 9'hdf == io_in_pc_bits[10:2] ? regs__223 : _GEN_225; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_227 = 9'he0 == io_in_pc_bits[10:2] ? regs__224 : _GEN_226; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_228 = 9'he1 == io_in_pc_bits[10:2] ? regs__225 : _GEN_227; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_229 = 9'he2 == io_in_pc_bits[10:2] ? regs__226 : _GEN_228; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_230 = 9'he3 == io_in_pc_bits[10:2] ? regs__227 : _GEN_229; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_231 = 9'he4 == io_in_pc_bits[10:2] ? regs__228 : _GEN_230; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_232 = 9'he5 == io_in_pc_bits[10:2] ? regs__229 : _GEN_231; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_233 = 9'he6 == io_in_pc_bits[10:2] ? regs__230 : _GEN_232; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_234 = 9'he7 == io_in_pc_bits[10:2] ? regs__231 : _GEN_233; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_235 = 9'he8 == io_in_pc_bits[10:2] ? regs__232 : _GEN_234; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_236 = 9'he9 == io_in_pc_bits[10:2] ? regs__233 : _GEN_235; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_237 = 9'hea == io_in_pc_bits[10:2] ? regs__234 : _GEN_236; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_238 = 9'heb == io_in_pc_bits[10:2] ? regs__235 : _GEN_237; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_239 = 9'hec == io_in_pc_bits[10:2] ? regs__236 : _GEN_238; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_240 = 9'hed == io_in_pc_bits[10:2] ? regs__237 : _GEN_239; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_241 = 9'hee == io_in_pc_bits[10:2] ? regs__238 : _GEN_240; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_242 = 9'hef == io_in_pc_bits[10:2] ? regs__239 : _GEN_241; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_243 = 9'hf0 == io_in_pc_bits[10:2] ? regs__240 : _GEN_242; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_244 = 9'hf1 == io_in_pc_bits[10:2] ? regs__241 : _GEN_243; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_245 = 9'hf2 == io_in_pc_bits[10:2] ? regs__242 : _GEN_244; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_246 = 9'hf3 == io_in_pc_bits[10:2] ? regs__243 : _GEN_245; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_247 = 9'hf4 == io_in_pc_bits[10:2] ? regs__244 : _GEN_246; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_248 = 9'hf5 == io_in_pc_bits[10:2] ? regs__245 : _GEN_247; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_249 = 9'hf6 == io_in_pc_bits[10:2] ? regs__246 : _GEN_248; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_250 = 9'hf7 == io_in_pc_bits[10:2] ? regs__247 : _GEN_249; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_251 = 9'hf8 == io_in_pc_bits[10:2] ? regs__248 : _GEN_250; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_252 = 9'hf9 == io_in_pc_bits[10:2] ? regs__249 : _GEN_251; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_253 = 9'hfa == io_in_pc_bits[10:2] ? regs__250 : _GEN_252; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_254 = 9'hfb == io_in_pc_bits[10:2] ? regs__251 : _GEN_253; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_255 = 9'hfc == io_in_pc_bits[10:2] ? regs__252 : _GEN_254; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_256 = 9'hfd == io_in_pc_bits[10:2] ? regs__253 : _GEN_255; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_257 = 9'hfe == io_in_pc_bits[10:2] ? regs__254 : _GEN_256; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_258 = 9'hff == io_in_pc_bits[10:2] ? regs__255 : _GEN_257; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_259 = 9'h100 == io_in_pc_bits[10:2] ? regs__256 : _GEN_258; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_260 = 9'h101 == io_in_pc_bits[10:2] ? regs__257 : _GEN_259; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_261 = 9'h102 == io_in_pc_bits[10:2] ? regs__258 : _GEN_260; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_262 = 9'h103 == io_in_pc_bits[10:2] ? regs__259 : _GEN_261; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_263 = 9'h104 == io_in_pc_bits[10:2] ? regs__260 : _GEN_262; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_264 = 9'h105 == io_in_pc_bits[10:2] ? regs__261 : _GEN_263; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_265 = 9'h106 == io_in_pc_bits[10:2] ? regs__262 : _GEN_264; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_266 = 9'h107 == io_in_pc_bits[10:2] ? regs__263 : _GEN_265; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_267 = 9'h108 == io_in_pc_bits[10:2] ? regs__264 : _GEN_266; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_268 = 9'h109 == io_in_pc_bits[10:2] ? regs__265 : _GEN_267; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_269 = 9'h10a == io_in_pc_bits[10:2] ? regs__266 : _GEN_268; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_270 = 9'h10b == io_in_pc_bits[10:2] ? regs__267 : _GEN_269; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_271 = 9'h10c == io_in_pc_bits[10:2] ? regs__268 : _GEN_270; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_272 = 9'h10d == io_in_pc_bits[10:2] ? regs__269 : _GEN_271; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_273 = 9'h10e == io_in_pc_bits[10:2] ? regs__270 : _GEN_272; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_274 = 9'h10f == io_in_pc_bits[10:2] ? regs__271 : _GEN_273; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_275 = 9'h110 == io_in_pc_bits[10:2] ? regs__272 : _GEN_274; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_276 = 9'h111 == io_in_pc_bits[10:2] ? regs__273 : _GEN_275; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_277 = 9'h112 == io_in_pc_bits[10:2] ? regs__274 : _GEN_276; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_278 = 9'h113 == io_in_pc_bits[10:2] ? regs__275 : _GEN_277; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_279 = 9'h114 == io_in_pc_bits[10:2] ? regs__276 : _GEN_278; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_280 = 9'h115 == io_in_pc_bits[10:2] ? regs__277 : _GEN_279; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_281 = 9'h116 == io_in_pc_bits[10:2] ? regs__278 : _GEN_280; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_282 = 9'h117 == io_in_pc_bits[10:2] ? regs__279 : _GEN_281; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_283 = 9'h118 == io_in_pc_bits[10:2] ? regs__280 : _GEN_282; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_284 = 9'h119 == io_in_pc_bits[10:2] ? regs__281 : _GEN_283; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_285 = 9'h11a == io_in_pc_bits[10:2] ? regs__282 : _GEN_284; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_286 = 9'h11b == io_in_pc_bits[10:2] ? regs__283 : _GEN_285; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_287 = 9'h11c == io_in_pc_bits[10:2] ? regs__284 : _GEN_286; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_288 = 9'h11d == io_in_pc_bits[10:2] ? regs__285 : _GEN_287; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_289 = 9'h11e == io_in_pc_bits[10:2] ? regs__286 : _GEN_288; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_290 = 9'h11f == io_in_pc_bits[10:2] ? regs__287 : _GEN_289; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_291 = 9'h120 == io_in_pc_bits[10:2] ? regs__288 : _GEN_290; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_292 = 9'h121 == io_in_pc_bits[10:2] ? regs__289 : _GEN_291; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_293 = 9'h122 == io_in_pc_bits[10:2] ? regs__290 : _GEN_292; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_294 = 9'h123 == io_in_pc_bits[10:2] ? regs__291 : _GEN_293; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_295 = 9'h124 == io_in_pc_bits[10:2] ? regs__292 : _GEN_294; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_296 = 9'h125 == io_in_pc_bits[10:2] ? regs__293 : _GEN_295; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_297 = 9'h126 == io_in_pc_bits[10:2] ? regs__294 : _GEN_296; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_298 = 9'h127 == io_in_pc_bits[10:2] ? regs__295 : _GEN_297; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_299 = 9'h128 == io_in_pc_bits[10:2] ? regs__296 : _GEN_298; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_300 = 9'h129 == io_in_pc_bits[10:2] ? regs__297 : _GEN_299; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_301 = 9'h12a == io_in_pc_bits[10:2] ? regs__298 : _GEN_300; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_302 = 9'h12b == io_in_pc_bits[10:2] ? regs__299 : _GEN_301; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_303 = 9'h12c == io_in_pc_bits[10:2] ? regs__300 : _GEN_302; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_304 = 9'h12d == io_in_pc_bits[10:2] ? regs__301 : _GEN_303; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_305 = 9'h12e == io_in_pc_bits[10:2] ? regs__302 : _GEN_304; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_306 = 9'h12f == io_in_pc_bits[10:2] ? regs__303 : _GEN_305; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_307 = 9'h130 == io_in_pc_bits[10:2] ? regs__304 : _GEN_306; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_308 = 9'h131 == io_in_pc_bits[10:2] ? regs__305 : _GEN_307; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_309 = 9'h132 == io_in_pc_bits[10:2] ? regs__306 : _GEN_308; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_310 = 9'h133 == io_in_pc_bits[10:2] ? regs__307 : _GEN_309; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_311 = 9'h134 == io_in_pc_bits[10:2] ? regs__308 : _GEN_310; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_312 = 9'h135 == io_in_pc_bits[10:2] ? regs__309 : _GEN_311; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_313 = 9'h136 == io_in_pc_bits[10:2] ? regs__310 : _GEN_312; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_314 = 9'h137 == io_in_pc_bits[10:2] ? regs__311 : _GEN_313; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_315 = 9'h138 == io_in_pc_bits[10:2] ? regs__312 : _GEN_314; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_316 = 9'h139 == io_in_pc_bits[10:2] ? regs__313 : _GEN_315; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_317 = 9'h13a == io_in_pc_bits[10:2] ? regs__314 : _GEN_316; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_318 = 9'h13b == io_in_pc_bits[10:2] ? regs__315 : _GEN_317; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_319 = 9'h13c == io_in_pc_bits[10:2] ? regs__316 : _GEN_318; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_320 = 9'h13d == io_in_pc_bits[10:2] ? regs__317 : _GEN_319; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_321 = 9'h13e == io_in_pc_bits[10:2] ? regs__318 : _GEN_320; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_322 = 9'h13f == io_in_pc_bits[10:2] ? regs__319 : _GEN_321; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_323 = 9'h140 == io_in_pc_bits[10:2] ? regs__320 : _GEN_322; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_324 = 9'h141 == io_in_pc_bits[10:2] ? regs__321 : _GEN_323; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_325 = 9'h142 == io_in_pc_bits[10:2] ? regs__322 : _GEN_324; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_326 = 9'h143 == io_in_pc_bits[10:2] ? regs__323 : _GEN_325; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_327 = 9'h144 == io_in_pc_bits[10:2] ? regs__324 : _GEN_326; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_328 = 9'h145 == io_in_pc_bits[10:2] ? regs__325 : _GEN_327; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_329 = 9'h146 == io_in_pc_bits[10:2] ? regs__326 : _GEN_328; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_330 = 9'h147 == io_in_pc_bits[10:2] ? regs__327 : _GEN_329; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_331 = 9'h148 == io_in_pc_bits[10:2] ? regs__328 : _GEN_330; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_332 = 9'h149 == io_in_pc_bits[10:2] ? regs__329 : _GEN_331; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_333 = 9'h14a == io_in_pc_bits[10:2] ? regs__330 : _GEN_332; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_334 = 9'h14b == io_in_pc_bits[10:2] ? regs__331 : _GEN_333; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_335 = 9'h14c == io_in_pc_bits[10:2] ? regs__332 : _GEN_334; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_336 = 9'h14d == io_in_pc_bits[10:2] ? regs__333 : _GEN_335; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_337 = 9'h14e == io_in_pc_bits[10:2] ? regs__334 : _GEN_336; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_338 = 9'h14f == io_in_pc_bits[10:2] ? regs__335 : _GEN_337; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_339 = 9'h150 == io_in_pc_bits[10:2] ? regs__336 : _GEN_338; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_340 = 9'h151 == io_in_pc_bits[10:2] ? regs__337 : _GEN_339; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_341 = 9'h152 == io_in_pc_bits[10:2] ? regs__338 : _GEN_340; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_342 = 9'h153 == io_in_pc_bits[10:2] ? regs__339 : _GEN_341; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_343 = 9'h154 == io_in_pc_bits[10:2] ? regs__340 : _GEN_342; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_344 = 9'h155 == io_in_pc_bits[10:2] ? regs__341 : _GEN_343; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_345 = 9'h156 == io_in_pc_bits[10:2] ? regs__342 : _GEN_344; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_346 = 9'h157 == io_in_pc_bits[10:2] ? regs__343 : _GEN_345; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_347 = 9'h158 == io_in_pc_bits[10:2] ? regs__344 : _GEN_346; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_348 = 9'h159 == io_in_pc_bits[10:2] ? regs__345 : _GEN_347; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_349 = 9'h15a == io_in_pc_bits[10:2] ? regs__346 : _GEN_348; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_350 = 9'h15b == io_in_pc_bits[10:2] ? regs__347 : _GEN_349; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_351 = 9'h15c == io_in_pc_bits[10:2] ? regs__348 : _GEN_350; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_352 = 9'h15d == io_in_pc_bits[10:2] ? regs__349 : _GEN_351; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_353 = 9'h15e == io_in_pc_bits[10:2] ? regs__350 : _GEN_352; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_354 = 9'h15f == io_in_pc_bits[10:2] ? regs__351 : _GEN_353; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_355 = 9'h160 == io_in_pc_bits[10:2] ? regs__352 : _GEN_354; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_356 = 9'h161 == io_in_pc_bits[10:2] ? regs__353 : _GEN_355; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_357 = 9'h162 == io_in_pc_bits[10:2] ? regs__354 : _GEN_356; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_358 = 9'h163 == io_in_pc_bits[10:2] ? regs__355 : _GEN_357; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_359 = 9'h164 == io_in_pc_bits[10:2] ? regs__356 : _GEN_358; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_360 = 9'h165 == io_in_pc_bits[10:2] ? regs__357 : _GEN_359; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_361 = 9'h166 == io_in_pc_bits[10:2] ? regs__358 : _GEN_360; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_362 = 9'h167 == io_in_pc_bits[10:2] ? regs__359 : _GEN_361; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_363 = 9'h168 == io_in_pc_bits[10:2] ? regs__360 : _GEN_362; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_364 = 9'h169 == io_in_pc_bits[10:2] ? regs__361 : _GEN_363; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_365 = 9'h16a == io_in_pc_bits[10:2] ? regs__362 : _GEN_364; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_366 = 9'h16b == io_in_pc_bits[10:2] ? regs__363 : _GEN_365; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_367 = 9'h16c == io_in_pc_bits[10:2] ? regs__364 : _GEN_366; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_368 = 9'h16d == io_in_pc_bits[10:2] ? regs__365 : _GEN_367; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_369 = 9'h16e == io_in_pc_bits[10:2] ? regs__366 : _GEN_368; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_370 = 9'h16f == io_in_pc_bits[10:2] ? regs__367 : _GEN_369; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_371 = 9'h170 == io_in_pc_bits[10:2] ? regs__368 : _GEN_370; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_372 = 9'h171 == io_in_pc_bits[10:2] ? regs__369 : _GEN_371; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_373 = 9'h172 == io_in_pc_bits[10:2] ? regs__370 : _GEN_372; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_374 = 9'h173 == io_in_pc_bits[10:2] ? regs__371 : _GEN_373; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_375 = 9'h174 == io_in_pc_bits[10:2] ? regs__372 : _GEN_374; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_376 = 9'h175 == io_in_pc_bits[10:2] ? regs__373 : _GEN_375; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_377 = 9'h176 == io_in_pc_bits[10:2] ? regs__374 : _GEN_376; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_378 = 9'h177 == io_in_pc_bits[10:2] ? regs__375 : _GEN_377; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_379 = 9'h178 == io_in_pc_bits[10:2] ? regs__376 : _GEN_378; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_380 = 9'h179 == io_in_pc_bits[10:2] ? regs__377 : _GEN_379; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_381 = 9'h17a == io_in_pc_bits[10:2] ? regs__378 : _GEN_380; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_382 = 9'h17b == io_in_pc_bits[10:2] ? regs__379 : _GEN_381; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_383 = 9'h17c == io_in_pc_bits[10:2] ? regs__380 : _GEN_382; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_384 = 9'h17d == io_in_pc_bits[10:2] ? regs__381 : _GEN_383; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_385 = 9'h17e == io_in_pc_bits[10:2] ? regs__382 : _GEN_384; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_386 = 9'h17f == io_in_pc_bits[10:2] ? regs__383 : _GEN_385; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_387 = 9'h180 == io_in_pc_bits[10:2] ? regs__384 : _GEN_386; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_388 = 9'h181 == io_in_pc_bits[10:2] ? regs__385 : _GEN_387; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_389 = 9'h182 == io_in_pc_bits[10:2] ? regs__386 : _GEN_388; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_390 = 9'h183 == io_in_pc_bits[10:2] ? regs__387 : _GEN_389; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_391 = 9'h184 == io_in_pc_bits[10:2] ? regs__388 : _GEN_390; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_392 = 9'h185 == io_in_pc_bits[10:2] ? regs__389 : _GEN_391; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_393 = 9'h186 == io_in_pc_bits[10:2] ? regs__390 : _GEN_392; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_394 = 9'h187 == io_in_pc_bits[10:2] ? regs__391 : _GEN_393; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_395 = 9'h188 == io_in_pc_bits[10:2] ? regs__392 : _GEN_394; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_396 = 9'h189 == io_in_pc_bits[10:2] ? regs__393 : _GEN_395; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_397 = 9'h18a == io_in_pc_bits[10:2] ? regs__394 : _GEN_396; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_398 = 9'h18b == io_in_pc_bits[10:2] ? regs__395 : _GEN_397; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_399 = 9'h18c == io_in_pc_bits[10:2] ? regs__396 : _GEN_398; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_400 = 9'h18d == io_in_pc_bits[10:2] ? regs__397 : _GEN_399; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_401 = 9'h18e == io_in_pc_bits[10:2] ? regs__398 : _GEN_400; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_402 = 9'h18f == io_in_pc_bits[10:2] ? regs__399 : _GEN_401; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_403 = 9'h190 == io_in_pc_bits[10:2] ? regs__400 : _GEN_402; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_404 = 9'h191 == io_in_pc_bits[10:2] ? regs__401 : _GEN_403; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_405 = 9'h192 == io_in_pc_bits[10:2] ? regs__402 : _GEN_404; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_406 = 9'h193 == io_in_pc_bits[10:2] ? regs__403 : _GEN_405; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_407 = 9'h194 == io_in_pc_bits[10:2] ? regs__404 : _GEN_406; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_408 = 9'h195 == io_in_pc_bits[10:2] ? regs__405 : _GEN_407; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_409 = 9'h196 == io_in_pc_bits[10:2] ? regs__406 : _GEN_408; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_410 = 9'h197 == io_in_pc_bits[10:2] ? regs__407 : _GEN_409; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_411 = 9'h198 == io_in_pc_bits[10:2] ? regs__408 : _GEN_410; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_412 = 9'h199 == io_in_pc_bits[10:2] ? regs__409 : _GEN_411; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_413 = 9'h19a == io_in_pc_bits[10:2] ? regs__410 : _GEN_412; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_414 = 9'h19b == io_in_pc_bits[10:2] ? regs__411 : _GEN_413; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_415 = 9'h19c == io_in_pc_bits[10:2] ? regs__412 : _GEN_414; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_416 = 9'h19d == io_in_pc_bits[10:2] ? regs__413 : _GEN_415; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_417 = 9'h19e == io_in_pc_bits[10:2] ? regs__414 : _GEN_416; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_418 = 9'h19f == io_in_pc_bits[10:2] ? regs__415 : _GEN_417; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_419 = 9'h1a0 == io_in_pc_bits[10:2] ? regs__416 : _GEN_418; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_420 = 9'h1a1 == io_in_pc_bits[10:2] ? regs__417 : _GEN_419; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_421 = 9'h1a2 == io_in_pc_bits[10:2] ? regs__418 : _GEN_420; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_422 = 9'h1a3 == io_in_pc_bits[10:2] ? regs__419 : _GEN_421; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_423 = 9'h1a4 == io_in_pc_bits[10:2] ? regs__420 : _GEN_422; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_424 = 9'h1a5 == io_in_pc_bits[10:2] ? regs__421 : _GEN_423; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_425 = 9'h1a6 == io_in_pc_bits[10:2] ? regs__422 : _GEN_424; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_426 = 9'h1a7 == io_in_pc_bits[10:2] ? regs__423 : _GEN_425; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_427 = 9'h1a8 == io_in_pc_bits[10:2] ? regs__424 : _GEN_426; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_428 = 9'h1a9 == io_in_pc_bits[10:2] ? regs__425 : _GEN_427; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_429 = 9'h1aa == io_in_pc_bits[10:2] ? regs__426 : _GEN_428; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_430 = 9'h1ab == io_in_pc_bits[10:2] ? regs__427 : _GEN_429; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_431 = 9'h1ac == io_in_pc_bits[10:2] ? regs__428 : _GEN_430; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_432 = 9'h1ad == io_in_pc_bits[10:2] ? regs__429 : _GEN_431; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_433 = 9'h1ae == io_in_pc_bits[10:2] ? regs__430 : _GEN_432; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_434 = 9'h1af == io_in_pc_bits[10:2] ? regs__431 : _GEN_433; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_435 = 9'h1b0 == io_in_pc_bits[10:2] ? regs__432 : _GEN_434; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_436 = 9'h1b1 == io_in_pc_bits[10:2] ? regs__433 : _GEN_435; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_437 = 9'h1b2 == io_in_pc_bits[10:2] ? regs__434 : _GEN_436; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_438 = 9'h1b3 == io_in_pc_bits[10:2] ? regs__435 : _GEN_437; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_439 = 9'h1b4 == io_in_pc_bits[10:2] ? regs__436 : _GEN_438; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_440 = 9'h1b5 == io_in_pc_bits[10:2] ? regs__437 : _GEN_439; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_441 = 9'h1b6 == io_in_pc_bits[10:2] ? regs__438 : _GEN_440; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_442 = 9'h1b7 == io_in_pc_bits[10:2] ? regs__439 : _GEN_441; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_443 = 9'h1b8 == io_in_pc_bits[10:2] ? regs__440 : _GEN_442; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_444 = 9'h1b9 == io_in_pc_bits[10:2] ? regs__441 : _GEN_443; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_445 = 9'h1ba == io_in_pc_bits[10:2] ? regs__442 : _GEN_444; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_446 = 9'h1bb == io_in_pc_bits[10:2] ? regs__443 : _GEN_445; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_447 = 9'h1bc == io_in_pc_bits[10:2] ? regs__444 : _GEN_446; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_448 = 9'h1bd == io_in_pc_bits[10:2] ? regs__445 : _GEN_447; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_449 = 9'h1be == io_in_pc_bits[10:2] ? regs__446 : _GEN_448; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_450 = 9'h1bf == io_in_pc_bits[10:2] ? regs__447 : _GEN_449; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_451 = 9'h1c0 == io_in_pc_bits[10:2] ? regs__448 : _GEN_450; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_452 = 9'h1c1 == io_in_pc_bits[10:2] ? regs__449 : _GEN_451; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_453 = 9'h1c2 == io_in_pc_bits[10:2] ? regs__450 : _GEN_452; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_454 = 9'h1c3 == io_in_pc_bits[10:2] ? regs__451 : _GEN_453; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_455 = 9'h1c4 == io_in_pc_bits[10:2] ? regs__452 : _GEN_454; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_456 = 9'h1c5 == io_in_pc_bits[10:2] ? regs__453 : _GEN_455; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_457 = 9'h1c6 == io_in_pc_bits[10:2] ? regs__454 : _GEN_456; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_458 = 9'h1c7 == io_in_pc_bits[10:2] ? regs__455 : _GEN_457; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_459 = 9'h1c8 == io_in_pc_bits[10:2] ? regs__456 : _GEN_458; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_460 = 9'h1c9 == io_in_pc_bits[10:2] ? regs__457 : _GEN_459; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_461 = 9'h1ca == io_in_pc_bits[10:2] ? regs__458 : _GEN_460; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_462 = 9'h1cb == io_in_pc_bits[10:2] ? regs__459 : _GEN_461; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_463 = 9'h1cc == io_in_pc_bits[10:2] ? regs__460 : _GEN_462; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_464 = 9'h1cd == io_in_pc_bits[10:2] ? regs__461 : _GEN_463; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_465 = 9'h1ce == io_in_pc_bits[10:2] ? regs__462 : _GEN_464; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_466 = 9'h1cf == io_in_pc_bits[10:2] ? regs__463 : _GEN_465; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_467 = 9'h1d0 == io_in_pc_bits[10:2] ? regs__464 : _GEN_466; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_468 = 9'h1d1 == io_in_pc_bits[10:2] ? regs__465 : _GEN_467; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_469 = 9'h1d2 == io_in_pc_bits[10:2] ? regs__466 : _GEN_468; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_470 = 9'h1d3 == io_in_pc_bits[10:2] ? regs__467 : _GEN_469; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_471 = 9'h1d4 == io_in_pc_bits[10:2] ? regs__468 : _GEN_470; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_472 = 9'h1d5 == io_in_pc_bits[10:2] ? regs__469 : _GEN_471; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_473 = 9'h1d6 == io_in_pc_bits[10:2] ? regs__470 : _GEN_472; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_474 = 9'h1d7 == io_in_pc_bits[10:2] ? regs__471 : _GEN_473; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_475 = 9'h1d8 == io_in_pc_bits[10:2] ? regs__472 : _GEN_474; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_476 = 9'h1d9 == io_in_pc_bits[10:2] ? regs__473 : _GEN_475; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_477 = 9'h1da == io_in_pc_bits[10:2] ? regs__474 : _GEN_476; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_478 = 9'h1db == io_in_pc_bits[10:2] ? regs__475 : _GEN_477; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_479 = 9'h1dc == io_in_pc_bits[10:2] ? regs__476 : _GEN_478; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_480 = 9'h1dd == io_in_pc_bits[10:2] ? regs__477 : _GEN_479; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_481 = 9'h1de == io_in_pc_bits[10:2] ? regs__478 : _GEN_480; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_482 = 9'h1df == io_in_pc_bits[10:2] ? regs__479 : _GEN_481; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_483 = 9'h1e0 == io_in_pc_bits[10:2] ? regs__480 : _GEN_482; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_484 = 9'h1e1 == io_in_pc_bits[10:2] ? regs__481 : _GEN_483; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_485 = 9'h1e2 == io_in_pc_bits[10:2] ? regs__482 : _GEN_484; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_486 = 9'h1e3 == io_in_pc_bits[10:2] ? regs__483 : _GEN_485; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_487 = 9'h1e4 == io_in_pc_bits[10:2] ? regs__484 : _GEN_486; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_488 = 9'h1e5 == io_in_pc_bits[10:2] ? regs__485 : _GEN_487; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_489 = 9'h1e6 == io_in_pc_bits[10:2] ? regs__486 : _GEN_488; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_490 = 9'h1e7 == io_in_pc_bits[10:2] ? regs__487 : _GEN_489; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_491 = 9'h1e8 == io_in_pc_bits[10:2] ? regs__488 : _GEN_490; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_492 = 9'h1e9 == io_in_pc_bits[10:2] ? regs__489 : _GEN_491; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_493 = 9'h1ea == io_in_pc_bits[10:2] ? regs__490 : _GEN_492; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_494 = 9'h1eb == io_in_pc_bits[10:2] ? regs__491 : _GEN_493; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_495 = 9'h1ec == io_in_pc_bits[10:2] ? regs__492 : _GEN_494; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_496 = 9'h1ed == io_in_pc_bits[10:2] ? regs__493 : _GEN_495; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_497 = 9'h1ee == io_in_pc_bits[10:2] ? regs__494 : _GEN_496; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_498 = 9'h1ef == io_in_pc_bits[10:2] ? regs__495 : _GEN_497; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_499 = 9'h1f0 == io_in_pc_bits[10:2] ? regs__496 : _GEN_498; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_500 = 9'h1f1 == io_in_pc_bits[10:2] ? regs__497 : _GEN_499; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_501 = 9'h1f2 == io_in_pc_bits[10:2] ? regs__498 : _GEN_500; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_502 = 9'h1f3 == io_in_pc_bits[10:2] ? regs__499 : _GEN_501; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_503 = 9'h1f4 == io_in_pc_bits[10:2] ? regs__500 : _GEN_502; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_504 = 9'h1f5 == io_in_pc_bits[10:2] ? regs__501 : _GEN_503; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_505 = 9'h1f6 == io_in_pc_bits[10:2] ? regs__502 : _GEN_504; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_506 = 9'h1f7 == io_in_pc_bits[10:2] ? regs__503 : _GEN_505; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_507 = 9'h1f8 == io_in_pc_bits[10:2] ? regs__504 : _GEN_506; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_508 = 9'h1f9 == io_in_pc_bits[10:2] ? regs__505 : _GEN_507; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_509 = 9'h1fa == io_in_pc_bits[10:2] ? regs__506 : _GEN_508; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_510 = 9'h1fb == io_in_pc_bits[10:2] ? regs__507 : _GEN_509; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_511 = 9'h1fc == io_in_pc_bits[10:2] ? regs__508 : _GEN_510; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_512 = 9'h1fd == io_in_pc_bits[10:2] ? regs__509 : _GEN_511; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_513 = 9'h1fe == io_in_pc_bits[10:2] ? regs__510 : _GEN_512; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  wire [1:0] _GEN_514 = 9'h1ff == io_in_pc_bits[10:2] ? regs__511 : _GEN_513; // @[src/main/scala/nutcore/frontend/BPU.scala 337:{67,67}]
  reg  phtTaken; // @[src/main/scala/nutcore/frontend/BPU.scala 337:27]
  reg [38:0] regs_1_0; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [38:0] regs_1_1; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [38:0] regs_1_2; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [38:0] regs_1_3; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [38:0] regs_1_4; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [38:0] regs_1_5; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [38:0] regs_1_6; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [38:0] regs_1_7; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [38:0] regs_1_8; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [38:0] regs_1_9; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [38:0] regs_1_10; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [38:0] regs_1_11; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [38:0] regs_1_12; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [38:0] regs_1_13; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [38:0] regs_1_14; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [38:0] regs_1_15; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [3:0] sp_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg [38:0] rasTarget; // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
  wire [38:0] _GEN_517 = 4'h1 == sp_value ? regs_1_1 : regs_1_0; // @[src/main/scala/nutcore/frontend/BPU.scala 345:{28,28}]
  wire [38:0] _GEN_518 = 4'h2 == sp_value ? regs_1_2 : _GEN_517; // @[src/main/scala/nutcore/frontend/BPU.scala 345:{28,28}]
  wire [38:0] _GEN_519 = 4'h3 == sp_value ? regs_1_3 : _GEN_518; // @[src/main/scala/nutcore/frontend/BPU.scala 345:{28,28}]
  wire [38:0] _GEN_520 = 4'h4 == sp_value ? regs_1_4 : _GEN_519; // @[src/main/scala/nutcore/frontend/BPU.scala 345:{28,28}]
  wire [38:0] _GEN_521 = 4'h5 == sp_value ? regs_1_5 : _GEN_520; // @[src/main/scala/nutcore/frontend/BPU.scala 345:{28,28}]
  wire [38:0] _GEN_522 = 4'h6 == sp_value ? regs_1_6 : _GEN_521; // @[src/main/scala/nutcore/frontend/BPU.scala 345:{28,28}]
  wire [38:0] _GEN_523 = 4'h7 == sp_value ? regs_1_7 : _GEN_522; // @[src/main/scala/nutcore/frontend/BPU.scala 345:{28,28}]
  wire [38:0] _GEN_524 = 4'h8 == sp_value ? regs_1_8 : _GEN_523; // @[src/main/scala/nutcore/frontend/BPU.scala 345:{28,28}]
  wire [38:0] _GEN_525 = 4'h9 == sp_value ? regs_1_9 : _GEN_524; // @[src/main/scala/nutcore/frontend/BPU.scala 345:{28,28}]
  wire [38:0] _GEN_526 = 4'ha == sp_value ? regs_1_10 : _GEN_525; // @[src/main/scala/nutcore/frontend/BPU.scala 345:{28,28}]
  wire [38:0] _GEN_527 = 4'hb == sp_value ? regs_1_11 : _GEN_526; // @[src/main/scala/nutcore/frontend/BPU.scala 345:{28,28}]
  wire [38:0] _GEN_528 = 4'hc == sp_value ? regs_1_12 : _GEN_527; // @[src/main/scala/nutcore/frontend/BPU.scala 345:{28,28}]
  wire  _T_35 = ~bpuUpdateReq_pc[1]; // @[src/main/scala/nutcore/frontend/BPU.scala 353:150]
  wire  _btbWrite_brIdx_T_3 = bpuUpdateReq_pc[2:0] == 3'h6 & ~bpuUpdateReq_isRVC; // @[src/main/scala/nutcore/frontend/BPU.scala 367:46]
  wire [1:0] btbWrite_brIdx_hi = {_btbWrite_brIdx_T_3,bpuUpdateReq_pc[1]}; // @[src/main/scala/nutcore/frontend/BPU.scala 367:24]
  reg [1:0] cnt; // @[src/main/scala/nutcore/frontend/BPU.scala 389:20]
  wire [1:0] _GEN_534 = 9'h1 == bpuUpdateReq_pc[10:2] ? regs__1 : regs__0; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_535 = 9'h2 == bpuUpdateReq_pc[10:2] ? regs__2 : _GEN_534; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_536 = 9'h3 == bpuUpdateReq_pc[10:2] ? regs__3 : _GEN_535; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_537 = 9'h4 == bpuUpdateReq_pc[10:2] ? regs__4 : _GEN_536; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_538 = 9'h5 == bpuUpdateReq_pc[10:2] ? regs__5 : _GEN_537; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_539 = 9'h6 == bpuUpdateReq_pc[10:2] ? regs__6 : _GEN_538; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_540 = 9'h7 == bpuUpdateReq_pc[10:2] ? regs__7 : _GEN_539; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_541 = 9'h8 == bpuUpdateReq_pc[10:2] ? regs__8 : _GEN_540; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_542 = 9'h9 == bpuUpdateReq_pc[10:2] ? regs__9 : _GEN_541; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_543 = 9'ha == bpuUpdateReq_pc[10:2] ? regs__10 : _GEN_542; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_544 = 9'hb == bpuUpdateReq_pc[10:2] ? regs__11 : _GEN_543; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_545 = 9'hc == bpuUpdateReq_pc[10:2] ? regs__12 : _GEN_544; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_546 = 9'hd == bpuUpdateReq_pc[10:2] ? regs__13 : _GEN_545; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_547 = 9'he == bpuUpdateReq_pc[10:2] ? regs__14 : _GEN_546; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_548 = 9'hf == bpuUpdateReq_pc[10:2] ? regs__15 : _GEN_547; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_549 = 9'h10 == bpuUpdateReq_pc[10:2] ? regs__16 : _GEN_548; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_550 = 9'h11 == bpuUpdateReq_pc[10:2] ? regs__17 : _GEN_549; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_551 = 9'h12 == bpuUpdateReq_pc[10:2] ? regs__18 : _GEN_550; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_552 = 9'h13 == bpuUpdateReq_pc[10:2] ? regs__19 : _GEN_551; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_553 = 9'h14 == bpuUpdateReq_pc[10:2] ? regs__20 : _GEN_552; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_554 = 9'h15 == bpuUpdateReq_pc[10:2] ? regs__21 : _GEN_553; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_555 = 9'h16 == bpuUpdateReq_pc[10:2] ? regs__22 : _GEN_554; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_556 = 9'h17 == bpuUpdateReq_pc[10:2] ? regs__23 : _GEN_555; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_557 = 9'h18 == bpuUpdateReq_pc[10:2] ? regs__24 : _GEN_556; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_558 = 9'h19 == bpuUpdateReq_pc[10:2] ? regs__25 : _GEN_557; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_559 = 9'h1a == bpuUpdateReq_pc[10:2] ? regs__26 : _GEN_558; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_560 = 9'h1b == bpuUpdateReq_pc[10:2] ? regs__27 : _GEN_559; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_561 = 9'h1c == bpuUpdateReq_pc[10:2] ? regs__28 : _GEN_560; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_562 = 9'h1d == bpuUpdateReq_pc[10:2] ? regs__29 : _GEN_561; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_563 = 9'h1e == bpuUpdateReq_pc[10:2] ? regs__30 : _GEN_562; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_564 = 9'h1f == bpuUpdateReq_pc[10:2] ? regs__31 : _GEN_563; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_565 = 9'h20 == bpuUpdateReq_pc[10:2] ? regs__32 : _GEN_564; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_566 = 9'h21 == bpuUpdateReq_pc[10:2] ? regs__33 : _GEN_565; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_567 = 9'h22 == bpuUpdateReq_pc[10:2] ? regs__34 : _GEN_566; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_568 = 9'h23 == bpuUpdateReq_pc[10:2] ? regs__35 : _GEN_567; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_569 = 9'h24 == bpuUpdateReq_pc[10:2] ? regs__36 : _GEN_568; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_570 = 9'h25 == bpuUpdateReq_pc[10:2] ? regs__37 : _GEN_569; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_571 = 9'h26 == bpuUpdateReq_pc[10:2] ? regs__38 : _GEN_570; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_572 = 9'h27 == bpuUpdateReq_pc[10:2] ? regs__39 : _GEN_571; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_573 = 9'h28 == bpuUpdateReq_pc[10:2] ? regs__40 : _GEN_572; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_574 = 9'h29 == bpuUpdateReq_pc[10:2] ? regs__41 : _GEN_573; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_575 = 9'h2a == bpuUpdateReq_pc[10:2] ? regs__42 : _GEN_574; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_576 = 9'h2b == bpuUpdateReq_pc[10:2] ? regs__43 : _GEN_575; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_577 = 9'h2c == bpuUpdateReq_pc[10:2] ? regs__44 : _GEN_576; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_578 = 9'h2d == bpuUpdateReq_pc[10:2] ? regs__45 : _GEN_577; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_579 = 9'h2e == bpuUpdateReq_pc[10:2] ? regs__46 : _GEN_578; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_580 = 9'h2f == bpuUpdateReq_pc[10:2] ? regs__47 : _GEN_579; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_581 = 9'h30 == bpuUpdateReq_pc[10:2] ? regs__48 : _GEN_580; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_582 = 9'h31 == bpuUpdateReq_pc[10:2] ? regs__49 : _GEN_581; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_583 = 9'h32 == bpuUpdateReq_pc[10:2] ? regs__50 : _GEN_582; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_584 = 9'h33 == bpuUpdateReq_pc[10:2] ? regs__51 : _GEN_583; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_585 = 9'h34 == bpuUpdateReq_pc[10:2] ? regs__52 : _GEN_584; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_586 = 9'h35 == bpuUpdateReq_pc[10:2] ? regs__53 : _GEN_585; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_587 = 9'h36 == bpuUpdateReq_pc[10:2] ? regs__54 : _GEN_586; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_588 = 9'h37 == bpuUpdateReq_pc[10:2] ? regs__55 : _GEN_587; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_589 = 9'h38 == bpuUpdateReq_pc[10:2] ? regs__56 : _GEN_588; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_590 = 9'h39 == bpuUpdateReq_pc[10:2] ? regs__57 : _GEN_589; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_591 = 9'h3a == bpuUpdateReq_pc[10:2] ? regs__58 : _GEN_590; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_592 = 9'h3b == bpuUpdateReq_pc[10:2] ? regs__59 : _GEN_591; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_593 = 9'h3c == bpuUpdateReq_pc[10:2] ? regs__60 : _GEN_592; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_594 = 9'h3d == bpuUpdateReq_pc[10:2] ? regs__61 : _GEN_593; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_595 = 9'h3e == bpuUpdateReq_pc[10:2] ? regs__62 : _GEN_594; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_596 = 9'h3f == bpuUpdateReq_pc[10:2] ? regs__63 : _GEN_595; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_597 = 9'h40 == bpuUpdateReq_pc[10:2] ? regs__64 : _GEN_596; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_598 = 9'h41 == bpuUpdateReq_pc[10:2] ? regs__65 : _GEN_597; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_599 = 9'h42 == bpuUpdateReq_pc[10:2] ? regs__66 : _GEN_598; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_600 = 9'h43 == bpuUpdateReq_pc[10:2] ? regs__67 : _GEN_599; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_601 = 9'h44 == bpuUpdateReq_pc[10:2] ? regs__68 : _GEN_600; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_602 = 9'h45 == bpuUpdateReq_pc[10:2] ? regs__69 : _GEN_601; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_603 = 9'h46 == bpuUpdateReq_pc[10:2] ? regs__70 : _GEN_602; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_604 = 9'h47 == bpuUpdateReq_pc[10:2] ? regs__71 : _GEN_603; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_605 = 9'h48 == bpuUpdateReq_pc[10:2] ? regs__72 : _GEN_604; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_606 = 9'h49 == bpuUpdateReq_pc[10:2] ? regs__73 : _GEN_605; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_607 = 9'h4a == bpuUpdateReq_pc[10:2] ? regs__74 : _GEN_606; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_608 = 9'h4b == bpuUpdateReq_pc[10:2] ? regs__75 : _GEN_607; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_609 = 9'h4c == bpuUpdateReq_pc[10:2] ? regs__76 : _GEN_608; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_610 = 9'h4d == bpuUpdateReq_pc[10:2] ? regs__77 : _GEN_609; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_611 = 9'h4e == bpuUpdateReq_pc[10:2] ? regs__78 : _GEN_610; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_612 = 9'h4f == bpuUpdateReq_pc[10:2] ? regs__79 : _GEN_611; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_613 = 9'h50 == bpuUpdateReq_pc[10:2] ? regs__80 : _GEN_612; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_614 = 9'h51 == bpuUpdateReq_pc[10:2] ? regs__81 : _GEN_613; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_615 = 9'h52 == bpuUpdateReq_pc[10:2] ? regs__82 : _GEN_614; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_616 = 9'h53 == bpuUpdateReq_pc[10:2] ? regs__83 : _GEN_615; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_617 = 9'h54 == bpuUpdateReq_pc[10:2] ? regs__84 : _GEN_616; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_618 = 9'h55 == bpuUpdateReq_pc[10:2] ? regs__85 : _GEN_617; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_619 = 9'h56 == bpuUpdateReq_pc[10:2] ? regs__86 : _GEN_618; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_620 = 9'h57 == bpuUpdateReq_pc[10:2] ? regs__87 : _GEN_619; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_621 = 9'h58 == bpuUpdateReq_pc[10:2] ? regs__88 : _GEN_620; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_622 = 9'h59 == bpuUpdateReq_pc[10:2] ? regs__89 : _GEN_621; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_623 = 9'h5a == bpuUpdateReq_pc[10:2] ? regs__90 : _GEN_622; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_624 = 9'h5b == bpuUpdateReq_pc[10:2] ? regs__91 : _GEN_623; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_625 = 9'h5c == bpuUpdateReq_pc[10:2] ? regs__92 : _GEN_624; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_626 = 9'h5d == bpuUpdateReq_pc[10:2] ? regs__93 : _GEN_625; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_627 = 9'h5e == bpuUpdateReq_pc[10:2] ? regs__94 : _GEN_626; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_628 = 9'h5f == bpuUpdateReq_pc[10:2] ? regs__95 : _GEN_627; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_629 = 9'h60 == bpuUpdateReq_pc[10:2] ? regs__96 : _GEN_628; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_630 = 9'h61 == bpuUpdateReq_pc[10:2] ? regs__97 : _GEN_629; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_631 = 9'h62 == bpuUpdateReq_pc[10:2] ? regs__98 : _GEN_630; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_632 = 9'h63 == bpuUpdateReq_pc[10:2] ? regs__99 : _GEN_631; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_633 = 9'h64 == bpuUpdateReq_pc[10:2] ? regs__100 : _GEN_632; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_634 = 9'h65 == bpuUpdateReq_pc[10:2] ? regs__101 : _GEN_633; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_635 = 9'h66 == bpuUpdateReq_pc[10:2] ? regs__102 : _GEN_634; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_636 = 9'h67 == bpuUpdateReq_pc[10:2] ? regs__103 : _GEN_635; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_637 = 9'h68 == bpuUpdateReq_pc[10:2] ? regs__104 : _GEN_636; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_638 = 9'h69 == bpuUpdateReq_pc[10:2] ? regs__105 : _GEN_637; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_639 = 9'h6a == bpuUpdateReq_pc[10:2] ? regs__106 : _GEN_638; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_640 = 9'h6b == bpuUpdateReq_pc[10:2] ? regs__107 : _GEN_639; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_641 = 9'h6c == bpuUpdateReq_pc[10:2] ? regs__108 : _GEN_640; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_642 = 9'h6d == bpuUpdateReq_pc[10:2] ? regs__109 : _GEN_641; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_643 = 9'h6e == bpuUpdateReq_pc[10:2] ? regs__110 : _GEN_642; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_644 = 9'h6f == bpuUpdateReq_pc[10:2] ? regs__111 : _GEN_643; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_645 = 9'h70 == bpuUpdateReq_pc[10:2] ? regs__112 : _GEN_644; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_646 = 9'h71 == bpuUpdateReq_pc[10:2] ? regs__113 : _GEN_645; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_647 = 9'h72 == bpuUpdateReq_pc[10:2] ? regs__114 : _GEN_646; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_648 = 9'h73 == bpuUpdateReq_pc[10:2] ? regs__115 : _GEN_647; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_649 = 9'h74 == bpuUpdateReq_pc[10:2] ? regs__116 : _GEN_648; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_650 = 9'h75 == bpuUpdateReq_pc[10:2] ? regs__117 : _GEN_649; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_651 = 9'h76 == bpuUpdateReq_pc[10:2] ? regs__118 : _GEN_650; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_652 = 9'h77 == bpuUpdateReq_pc[10:2] ? regs__119 : _GEN_651; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_653 = 9'h78 == bpuUpdateReq_pc[10:2] ? regs__120 : _GEN_652; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_654 = 9'h79 == bpuUpdateReq_pc[10:2] ? regs__121 : _GEN_653; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_655 = 9'h7a == bpuUpdateReq_pc[10:2] ? regs__122 : _GEN_654; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_656 = 9'h7b == bpuUpdateReq_pc[10:2] ? regs__123 : _GEN_655; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_657 = 9'h7c == bpuUpdateReq_pc[10:2] ? regs__124 : _GEN_656; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_658 = 9'h7d == bpuUpdateReq_pc[10:2] ? regs__125 : _GEN_657; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_659 = 9'h7e == bpuUpdateReq_pc[10:2] ? regs__126 : _GEN_658; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_660 = 9'h7f == bpuUpdateReq_pc[10:2] ? regs__127 : _GEN_659; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_661 = 9'h80 == bpuUpdateReq_pc[10:2] ? regs__128 : _GEN_660; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_662 = 9'h81 == bpuUpdateReq_pc[10:2] ? regs__129 : _GEN_661; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_663 = 9'h82 == bpuUpdateReq_pc[10:2] ? regs__130 : _GEN_662; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_664 = 9'h83 == bpuUpdateReq_pc[10:2] ? regs__131 : _GEN_663; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_665 = 9'h84 == bpuUpdateReq_pc[10:2] ? regs__132 : _GEN_664; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_666 = 9'h85 == bpuUpdateReq_pc[10:2] ? regs__133 : _GEN_665; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_667 = 9'h86 == bpuUpdateReq_pc[10:2] ? regs__134 : _GEN_666; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_668 = 9'h87 == bpuUpdateReq_pc[10:2] ? regs__135 : _GEN_667; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_669 = 9'h88 == bpuUpdateReq_pc[10:2] ? regs__136 : _GEN_668; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_670 = 9'h89 == bpuUpdateReq_pc[10:2] ? regs__137 : _GEN_669; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_671 = 9'h8a == bpuUpdateReq_pc[10:2] ? regs__138 : _GEN_670; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_672 = 9'h8b == bpuUpdateReq_pc[10:2] ? regs__139 : _GEN_671; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_673 = 9'h8c == bpuUpdateReq_pc[10:2] ? regs__140 : _GEN_672; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_674 = 9'h8d == bpuUpdateReq_pc[10:2] ? regs__141 : _GEN_673; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_675 = 9'h8e == bpuUpdateReq_pc[10:2] ? regs__142 : _GEN_674; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_676 = 9'h8f == bpuUpdateReq_pc[10:2] ? regs__143 : _GEN_675; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_677 = 9'h90 == bpuUpdateReq_pc[10:2] ? regs__144 : _GEN_676; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_678 = 9'h91 == bpuUpdateReq_pc[10:2] ? regs__145 : _GEN_677; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_679 = 9'h92 == bpuUpdateReq_pc[10:2] ? regs__146 : _GEN_678; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_680 = 9'h93 == bpuUpdateReq_pc[10:2] ? regs__147 : _GEN_679; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_681 = 9'h94 == bpuUpdateReq_pc[10:2] ? regs__148 : _GEN_680; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_682 = 9'h95 == bpuUpdateReq_pc[10:2] ? regs__149 : _GEN_681; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_683 = 9'h96 == bpuUpdateReq_pc[10:2] ? regs__150 : _GEN_682; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_684 = 9'h97 == bpuUpdateReq_pc[10:2] ? regs__151 : _GEN_683; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_685 = 9'h98 == bpuUpdateReq_pc[10:2] ? regs__152 : _GEN_684; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_686 = 9'h99 == bpuUpdateReq_pc[10:2] ? regs__153 : _GEN_685; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_687 = 9'h9a == bpuUpdateReq_pc[10:2] ? regs__154 : _GEN_686; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_688 = 9'h9b == bpuUpdateReq_pc[10:2] ? regs__155 : _GEN_687; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_689 = 9'h9c == bpuUpdateReq_pc[10:2] ? regs__156 : _GEN_688; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_690 = 9'h9d == bpuUpdateReq_pc[10:2] ? regs__157 : _GEN_689; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_691 = 9'h9e == bpuUpdateReq_pc[10:2] ? regs__158 : _GEN_690; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_692 = 9'h9f == bpuUpdateReq_pc[10:2] ? regs__159 : _GEN_691; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_693 = 9'ha0 == bpuUpdateReq_pc[10:2] ? regs__160 : _GEN_692; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_694 = 9'ha1 == bpuUpdateReq_pc[10:2] ? regs__161 : _GEN_693; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_695 = 9'ha2 == bpuUpdateReq_pc[10:2] ? regs__162 : _GEN_694; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_696 = 9'ha3 == bpuUpdateReq_pc[10:2] ? regs__163 : _GEN_695; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_697 = 9'ha4 == bpuUpdateReq_pc[10:2] ? regs__164 : _GEN_696; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_698 = 9'ha5 == bpuUpdateReq_pc[10:2] ? regs__165 : _GEN_697; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_699 = 9'ha6 == bpuUpdateReq_pc[10:2] ? regs__166 : _GEN_698; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_700 = 9'ha7 == bpuUpdateReq_pc[10:2] ? regs__167 : _GEN_699; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_701 = 9'ha8 == bpuUpdateReq_pc[10:2] ? regs__168 : _GEN_700; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_702 = 9'ha9 == bpuUpdateReq_pc[10:2] ? regs__169 : _GEN_701; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_703 = 9'haa == bpuUpdateReq_pc[10:2] ? regs__170 : _GEN_702; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_704 = 9'hab == bpuUpdateReq_pc[10:2] ? regs__171 : _GEN_703; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_705 = 9'hac == bpuUpdateReq_pc[10:2] ? regs__172 : _GEN_704; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_706 = 9'had == bpuUpdateReq_pc[10:2] ? regs__173 : _GEN_705; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_707 = 9'hae == bpuUpdateReq_pc[10:2] ? regs__174 : _GEN_706; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_708 = 9'haf == bpuUpdateReq_pc[10:2] ? regs__175 : _GEN_707; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_709 = 9'hb0 == bpuUpdateReq_pc[10:2] ? regs__176 : _GEN_708; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_710 = 9'hb1 == bpuUpdateReq_pc[10:2] ? regs__177 : _GEN_709; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_711 = 9'hb2 == bpuUpdateReq_pc[10:2] ? regs__178 : _GEN_710; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_712 = 9'hb3 == bpuUpdateReq_pc[10:2] ? regs__179 : _GEN_711; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_713 = 9'hb4 == bpuUpdateReq_pc[10:2] ? regs__180 : _GEN_712; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_714 = 9'hb5 == bpuUpdateReq_pc[10:2] ? regs__181 : _GEN_713; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_715 = 9'hb6 == bpuUpdateReq_pc[10:2] ? regs__182 : _GEN_714; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_716 = 9'hb7 == bpuUpdateReq_pc[10:2] ? regs__183 : _GEN_715; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_717 = 9'hb8 == bpuUpdateReq_pc[10:2] ? regs__184 : _GEN_716; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_718 = 9'hb9 == bpuUpdateReq_pc[10:2] ? regs__185 : _GEN_717; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_719 = 9'hba == bpuUpdateReq_pc[10:2] ? regs__186 : _GEN_718; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_720 = 9'hbb == bpuUpdateReq_pc[10:2] ? regs__187 : _GEN_719; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_721 = 9'hbc == bpuUpdateReq_pc[10:2] ? regs__188 : _GEN_720; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_722 = 9'hbd == bpuUpdateReq_pc[10:2] ? regs__189 : _GEN_721; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_723 = 9'hbe == bpuUpdateReq_pc[10:2] ? regs__190 : _GEN_722; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_724 = 9'hbf == bpuUpdateReq_pc[10:2] ? regs__191 : _GEN_723; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_725 = 9'hc0 == bpuUpdateReq_pc[10:2] ? regs__192 : _GEN_724; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_726 = 9'hc1 == bpuUpdateReq_pc[10:2] ? regs__193 : _GEN_725; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_727 = 9'hc2 == bpuUpdateReq_pc[10:2] ? regs__194 : _GEN_726; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_728 = 9'hc3 == bpuUpdateReq_pc[10:2] ? regs__195 : _GEN_727; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_729 = 9'hc4 == bpuUpdateReq_pc[10:2] ? regs__196 : _GEN_728; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_730 = 9'hc5 == bpuUpdateReq_pc[10:2] ? regs__197 : _GEN_729; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_731 = 9'hc6 == bpuUpdateReq_pc[10:2] ? regs__198 : _GEN_730; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_732 = 9'hc7 == bpuUpdateReq_pc[10:2] ? regs__199 : _GEN_731; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_733 = 9'hc8 == bpuUpdateReq_pc[10:2] ? regs__200 : _GEN_732; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_734 = 9'hc9 == bpuUpdateReq_pc[10:2] ? regs__201 : _GEN_733; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_735 = 9'hca == bpuUpdateReq_pc[10:2] ? regs__202 : _GEN_734; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_736 = 9'hcb == bpuUpdateReq_pc[10:2] ? regs__203 : _GEN_735; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_737 = 9'hcc == bpuUpdateReq_pc[10:2] ? regs__204 : _GEN_736; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_738 = 9'hcd == bpuUpdateReq_pc[10:2] ? regs__205 : _GEN_737; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_739 = 9'hce == bpuUpdateReq_pc[10:2] ? regs__206 : _GEN_738; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_740 = 9'hcf == bpuUpdateReq_pc[10:2] ? regs__207 : _GEN_739; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_741 = 9'hd0 == bpuUpdateReq_pc[10:2] ? regs__208 : _GEN_740; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_742 = 9'hd1 == bpuUpdateReq_pc[10:2] ? regs__209 : _GEN_741; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_743 = 9'hd2 == bpuUpdateReq_pc[10:2] ? regs__210 : _GEN_742; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_744 = 9'hd3 == bpuUpdateReq_pc[10:2] ? regs__211 : _GEN_743; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_745 = 9'hd4 == bpuUpdateReq_pc[10:2] ? regs__212 : _GEN_744; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_746 = 9'hd5 == bpuUpdateReq_pc[10:2] ? regs__213 : _GEN_745; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_747 = 9'hd6 == bpuUpdateReq_pc[10:2] ? regs__214 : _GEN_746; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_748 = 9'hd7 == bpuUpdateReq_pc[10:2] ? regs__215 : _GEN_747; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_749 = 9'hd8 == bpuUpdateReq_pc[10:2] ? regs__216 : _GEN_748; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_750 = 9'hd9 == bpuUpdateReq_pc[10:2] ? regs__217 : _GEN_749; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_751 = 9'hda == bpuUpdateReq_pc[10:2] ? regs__218 : _GEN_750; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_752 = 9'hdb == bpuUpdateReq_pc[10:2] ? regs__219 : _GEN_751; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_753 = 9'hdc == bpuUpdateReq_pc[10:2] ? regs__220 : _GEN_752; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_754 = 9'hdd == bpuUpdateReq_pc[10:2] ? regs__221 : _GEN_753; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_755 = 9'hde == bpuUpdateReq_pc[10:2] ? regs__222 : _GEN_754; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_756 = 9'hdf == bpuUpdateReq_pc[10:2] ? regs__223 : _GEN_755; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_757 = 9'he0 == bpuUpdateReq_pc[10:2] ? regs__224 : _GEN_756; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_758 = 9'he1 == bpuUpdateReq_pc[10:2] ? regs__225 : _GEN_757; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_759 = 9'he2 == bpuUpdateReq_pc[10:2] ? regs__226 : _GEN_758; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_760 = 9'he3 == bpuUpdateReq_pc[10:2] ? regs__227 : _GEN_759; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_761 = 9'he4 == bpuUpdateReq_pc[10:2] ? regs__228 : _GEN_760; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_762 = 9'he5 == bpuUpdateReq_pc[10:2] ? regs__229 : _GEN_761; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_763 = 9'he6 == bpuUpdateReq_pc[10:2] ? regs__230 : _GEN_762; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_764 = 9'he7 == bpuUpdateReq_pc[10:2] ? regs__231 : _GEN_763; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_765 = 9'he8 == bpuUpdateReq_pc[10:2] ? regs__232 : _GEN_764; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_766 = 9'he9 == bpuUpdateReq_pc[10:2] ? regs__233 : _GEN_765; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_767 = 9'hea == bpuUpdateReq_pc[10:2] ? regs__234 : _GEN_766; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_768 = 9'heb == bpuUpdateReq_pc[10:2] ? regs__235 : _GEN_767; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_769 = 9'hec == bpuUpdateReq_pc[10:2] ? regs__236 : _GEN_768; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_770 = 9'hed == bpuUpdateReq_pc[10:2] ? regs__237 : _GEN_769; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_771 = 9'hee == bpuUpdateReq_pc[10:2] ? regs__238 : _GEN_770; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_772 = 9'hef == bpuUpdateReq_pc[10:2] ? regs__239 : _GEN_771; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_773 = 9'hf0 == bpuUpdateReq_pc[10:2] ? regs__240 : _GEN_772; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_774 = 9'hf1 == bpuUpdateReq_pc[10:2] ? regs__241 : _GEN_773; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_775 = 9'hf2 == bpuUpdateReq_pc[10:2] ? regs__242 : _GEN_774; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_776 = 9'hf3 == bpuUpdateReq_pc[10:2] ? regs__243 : _GEN_775; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_777 = 9'hf4 == bpuUpdateReq_pc[10:2] ? regs__244 : _GEN_776; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_778 = 9'hf5 == bpuUpdateReq_pc[10:2] ? regs__245 : _GEN_777; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_779 = 9'hf6 == bpuUpdateReq_pc[10:2] ? regs__246 : _GEN_778; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_780 = 9'hf7 == bpuUpdateReq_pc[10:2] ? regs__247 : _GEN_779; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_781 = 9'hf8 == bpuUpdateReq_pc[10:2] ? regs__248 : _GEN_780; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_782 = 9'hf9 == bpuUpdateReq_pc[10:2] ? regs__249 : _GEN_781; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_783 = 9'hfa == bpuUpdateReq_pc[10:2] ? regs__250 : _GEN_782; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_784 = 9'hfb == bpuUpdateReq_pc[10:2] ? regs__251 : _GEN_783; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_785 = 9'hfc == bpuUpdateReq_pc[10:2] ? regs__252 : _GEN_784; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_786 = 9'hfd == bpuUpdateReq_pc[10:2] ? regs__253 : _GEN_785; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_787 = 9'hfe == bpuUpdateReq_pc[10:2] ? regs__254 : _GEN_786; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_788 = 9'hff == bpuUpdateReq_pc[10:2] ? regs__255 : _GEN_787; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_789 = 9'h100 == bpuUpdateReq_pc[10:2] ? regs__256 : _GEN_788; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_790 = 9'h101 == bpuUpdateReq_pc[10:2] ? regs__257 : _GEN_789; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_791 = 9'h102 == bpuUpdateReq_pc[10:2] ? regs__258 : _GEN_790; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_792 = 9'h103 == bpuUpdateReq_pc[10:2] ? regs__259 : _GEN_791; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_793 = 9'h104 == bpuUpdateReq_pc[10:2] ? regs__260 : _GEN_792; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_794 = 9'h105 == bpuUpdateReq_pc[10:2] ? regs__261 : _GEN_793; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_795 = 9'h106 == bpuUpdateReq_pc[10:2] ? regs__262 : _GEN_794; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_796 = 9'h107 == bpuUpdateReq_pc[10:2] ? regs__263 : _GEN_795; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_797 = 9'h108 == bpuUpdateReq_pc[10:2] ? regs__264 : _GEN_796; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_798 = 9'h109 == bpuUpdateReq_pc[10:2] ? regs__265 : _GEN_797; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_799 = 9'h10a == bpuUpdateReq_pc[10:2] ? regs__266 : _GEN_798; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_800 = 9'h10b == bpuUpdateReq_pc[10:2] ? regs__267 : _GEN_799; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_801 = 9'h10c == bpuUpdateReq_pc[10:2] ? regs__268 : _GEN_800; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_802 = 9'h10d == bpuUpdateReq_pc[10:2] ? regs__269 : _GEN_801; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_803 = 9'h10e == bpuUpdateReq_pc[10:2] ? regs__270 : _GEN_802; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_804 = 9'h10f == bpuUpdateReq_pc[10:2] ? regs__271 : _GEN_803; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_805 = 9'h110 == bpuUpdateReq_pc[10:2] ? regs__272 : _GEN_804; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_806 = 9'h111 == bpuUpdateReq_pc[10:2] ? regs__273 : _GEN_805; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_807 = 9'h112 == bpuUpdateReq_pc[10:2] ? regs__274 : _GEN_806; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_808 = 9'h113 == bpuUpdateReq_pc[10:2] ? regs__275 : _GEN_807; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_809 = 9'h114 == bpuUpdateReq_pc[10:2] ? regs__276 : _GEN_808; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_810 = 9'h115 == bpuUpdateReq_pc[10:2] ? regs__277 : _GEN_809; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_811 = 9'h116 == bpuUpdateReq_pc[10:2] ? regs__278 : _GEN_810; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_812 = 9'h117 == bpuUpdateReq_pc[10:2] ? regs__279 : _GEN_811; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_813 = 9'h118 == bpuUpdateReq_pc[10:2] ? regs__280 : _GEN_812; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_814 = 9'h119 == bpuUpdateReq_pc[10:2] ? regs__281 : _GEN_813; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_815 = 9'h11a == bpuUpdateReq_pc[10:2] ? regs__282 : _GEN_814; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_816 = 9'h11b == bpuUpdateReq_pc[10:2] ? regs__283 : _GEN_815; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_817 = 9'h11c == bpuUpdateReq_pc[10:2] ? regs__284 : _GEN_816; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_818 = 9'h11d == bpuUpdateReq_pc[10:2] ? regs__285 : _GEN_817; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_819 = 9'h11e == bpuUpdateReq_pc[10:2] ? regs__286 : _GEN_818; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_820 = 9'h11f == bpuUpdateReq_pc[10:2] ? regs__287 : _GEN_819; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_821 = 9'h120 == bpuUpdateReq_pc[10:2] ? regs__288 : _GEN_820; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_822 = 9'h121 == bpuUpdateReq_pc[10:2] ? regs__289 : _GEN_821; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_823 = 9'h122 == bpuUpdateReq_pc[10:2] ? regs__290 : _GEN_822; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_824 = 9'h123 == bpuUpdateReq_pc[10:2] ? regs__291 : _GEN_823; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_825 = 9'h124 == bpuUpdateReq_pc[10:2] ? regs__292 : _GEN_824; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_826 = 9'h125 == bpuUpdateReq_pc[10:2] ? regs__293 : _GEN_825; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_827 = 9'h126 == bpuUpdateReq_pc[10:2] ? regs__294 : _GEN_826; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_828 = 9'h127 == bpuUpdateReq_pc[10:2] ? regs__295 : _GEN_827; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_829 = 9'h128 == bpuUpdateReq_pc[10:2] ? regs__296 : _GEN_828; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_830 = 9'h129 == bpuUpdateReq_pc[10:2] ? regs__297 : _GEN_829; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_831 = 9'h12a == bpuUpdateReq_pc[10:2] ? regs__298 : _GEN_830; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_832 = 9'h12b == bpuUpdateReq_pc[10:2] ? regs__299 : _GEN_831; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_833 = 9'h12c == bpuUpdateReq_pc[10:2] ? regs__300 : _GEN_832; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_834 = 9'h12d == bpuUpdateReq_pc[10:2] ? regs__301 : _GEN_833; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_835 = 9'h12e == bpuUpdateReq_pc[10:2] ? regs__302 : _GEN_834; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_836 = 9'h12f == bpuUpdateReq_pc[10:2] ? regs__303 : _GEN_835; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_837 = 9'h130 == bpuUpdateReq_pc[10:2] ? regs__304 : _GEN_836; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_838 = 9'h131 == bpuUpdateReq_pc[10:2] ? regs__305 : _GEN_837; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_839 = 9'h132 == bpuUpdateReq_pc[10:2] ? regs__306 : _GEN_838; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_840 = 9'h133 == bpuUpdateReq_pc[10:2] ? regs__307 : _GEN_839; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_841 = 9'h134 == bpuUpdateReq_pc[10:2] ? regs__308 : _GEN_840; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_842 = 9'h135 == bpuUpdateReq_pc[10:2] ? regs__309 : _GEN_841; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_843 = 9'h136 == bpuUpdateReq_pc[10:2] ? regs__310 : _GEN_842; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_844 = 9'h137 == bpuUpdateReq_pc[10:2] ? regs__311 : _GEN_843; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_845 = 9'h138 == bpuUpdateReq_pc[10:2] ? regs__312 : _GEN_844; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_846 = 9'h139 == bpuUpdateReq_pc[10:2] ? regs__313 : _GEN_845; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_847 = 9'h13a == bpuUpdateReq_pc[10:2] ? regs__314 : _GEN_846; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_848 = 9'h13b == bpuUpdateReq_pc[10:2] ? regs__315 : _GEN_847; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_849 = 9'h13c == bpuUpdateReq_pc[10:2] ? regs__316 : _GEN_848; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_850 = 9'h13d == bpuUpdateReq_pc[10:2] ? regs__317 : _GEN_849; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_851 = 9'h13e == bpuUpdateReq_pc[10:2] ? regs__318 : _GEN_850; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_852 = 9'h13f == bpuUpdateReq_pc[10:2] ? regs__319 : _GEN_851; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_853 = 9'h140 == bpuUpdateReq_pc[10:2] ? regs__320 : _GEN_852; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_854 = 9'h141 == bpuUpdateReq_pc[10:2] ? regs__321 : _GEN_853; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_855 = 9'h142 == bpuUpdateReq_pc[10:2] ? regs__322 : _GEN_854; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_856 = 9'h143 == bpuUpdateReq_pc[10:2] ? regs__323 : _GEN_855; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_857 = 9'h144 == bpuUpdateReq_pc[10:2] ? regs__324 : _GEN_856; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_858 = 9'h145 == bpuUpdateReq_pc[10:2] ? regs__325 : _GEN_857; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_859 = 9'h146 == bpuUpdateReq_pc[10:2] ? regs__326 : _GEN_858; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_860 = 9'h147 == bpuUpdateReq_pc[10:2] ? regs__327 : _GEN_859; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_861 = 9'h148 == bpuUpdateReq_pc[10:2] ? regs__328 : _GEN_860; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_862 = 9'h149 == bpuUpdateReq_pc[10:2] ? regs__329 : _GEN_861; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_863 = 9'h14a == bpuUpdateReq_pc[10:2] ? regs__330 : _GEN_862; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_864 = 9'h14b == bpuUpdateReq_pc[10:2] ? regs__331 : _GEN_863; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_865 = 9'h14c == bpuUpdateReq_pc[10:2] ? regs__332 : _GEN_864; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_866 = 9'h14d == bpuUpdateReq_pc[10:2] ? regs__333 : _GEN_865; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_867 = 9'h14e == bpuUpdateReq_pc[10:2] ? regs__334 : _GEN_866; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_868 = 9'h14f == bpuUpdateReq_pc[10:2] ? regs__335 : _GEN_867; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_869 = 9'h150 == bpuUpdateReq_pc[10:2] ? regs__336 : _GEN_868; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_870 = 9'h151 == bpuUpdateReq_pc[10:2] ? regs__337 : _GEN_869; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_871 = 9'h152 == bpuUpdateReq_pc[10:2] ? regs__338 : _GEN_870; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_872 = 9'h153 == bpuUpdateReq_pc[10:2] ? regs__339 : _GEN_871; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_873 = 9'h154 == bpuUpdateReq_pc[10:2] ? regs__340 : _GEN_872; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_874 = 9'h155 == bpuUpdateReq_pc[10:2] ? regs__341 : _GEN_873; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_875 = 9'h156 == bpuUpdateReq_pc[10:2] ? regs__342 : _GEN_874; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_876 = 9'h157 == bpuUpdateReq_pc[10:2] ? regs__343 : _GEN_875; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_877 = 9'h158 == bpuUpdateReq_pc[10:2] ? regs__344 : _GEN_876; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_878 = 9'h159 == bpuUpdateReq_pc[10:2] ? regs__345 : _GEN_877; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_879 = 9'h15a == bpuUpdateReq_pc[10:2] ? regs__346 : _GEN_878; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_880 = 9'h15b == bpuUpdateReq_pc[10:2] ? regs__347 : _GEN_879; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_881 = 9'h15c == bpuUpdateReq_pc[10:2] ? regs__348 : _GEN_880; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_882 = 9'h15d == bpuUpdateReq_pc[10:2] ? regs__349 : _GEN_881; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_883 = 9'h15e == bpuUpdateReq_pc[10:2] ? regs__350 : _GEN_882; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_884 = 9'h15f == bpuUpdateReq_pc[10:2] ? regs__351 : _GEN_883; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_885 = 9'h160 == bpuUpdateReq_pc[10:2] ? regs__352 : _GEN_884; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_886 = 9'h161 == bpuUpdateReq_pc[10:2] ? regs__353 : _GEN_885; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_887 = 9'h162 == bpuUpdateReq_pc[10:2] ? regs__354 : _GEN_886; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_888 = 9'h163 == bpuUpdateReq_pc[10:2] ? regs__355 : _GEN_887; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_889 = 9'h164 == bpuUpdateReq_pc[10:2] ? regs__356 : _GEN_888; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_890 = 9'h165 == bpuUpdateReq_pc[10:2] ? regs__357 : _GEN_889; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_891 = 9'h166 == bpuUpdateReq_pc[10:2] ? regs__358 : _GEN_890; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_892 = 9'h167 == bpuUpdateReq_pc[10:2] ? regs__359 : _GEN_891; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_893 = 9'h168 == bpuUpdateReq_pc[10:2] ? regs__360 : _GEN_892; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_894 = 9'h169 == bpuUpdateReq_pc[10:2] ? regs__361 : _GEN_893; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_895 = 9'h16a == bpuUpdateReq_pc[10:2] ? regs__362 : _GEN_894; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_896 = 9'h16b == bpuUpdateReq_pc[10:2] ? regs__363 : _GEN_895; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_897 = 9'h16c == bpuUpdateReq_pc[10:2] ? regs__364 : _GEN_896; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_898 = 9'h16d == bpuUpdateReq_pc[10:2] ? regs__365 : _GEN_897; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_899 = 9'h16e == bpuUpdateReq_pc[10:2] ? regs__366 : _GEN_898; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_900 = 9'h16f == bpuUpdateReq_pc[10:2] ? regs__367 : _GEN_899; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_901 = 9'h170 == bpuUpdateReq_pc[10:2] ? regs__368 : _GEN_900; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_902 = 9'h171 == bpuUpdateReq_pc[10:2] ? regs__369 : _GEN_901; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_903 = 9'h172 == bpuUpdateReq_pc[10:2] ? regs__370 : _GEN_902; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_904 = 9'h173 == bpuUpdateReq_pc[10:2] ? regs__371 : _GEN_903; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_905 = 9'h174 == bpuUpdateReq_pc[10:2] ? regs__372 : _GEN_904; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_906 = 9'h175 == bpuUpdateReq_pc[10:2] ? regs__373 : _GEN_905; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_907 = 9'h176 == bpuUpdateReq_pc[10:2] ? regs__374 : _GEN_906; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_908 = 9'h177 == bpuUpdateReq_pc[10:2] ? regs__375 : _GEN_907; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_909 = 9'h178 == bpuUpdateReq_pc[10:2] ? regs__376 : _GEN_908; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_910 = 9'h179 == bpuUpdateReq_pc[10:2] ? regs__377 : _GEN_909; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_911 = 9'h17a == bpuUpdateReq_pc[10:2] ? regs__378 : _GEN_910; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_912 = 9'h17b == bpuUpdateReq_pc[10:2] ? regs__379 : _GEN_911; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_913 = 9'h17c == bpuUpdateReq_pc[10:2] ? regs__380 : _GEN_912; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_914 = 9'h17d == bpuUpdateReq_pc[10:2] ? regs__381 : _GEN_913; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_915 = 9'h17e == bpuUpdateReq_pc[10:2] ? regs__382 : _GEN_914; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_916 = 9'h17f == bpuUpdateReq_pc[10:2] ? regs__383 : _GEN_915; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_917 = 9'h180 == bpuUpdateReq_pc[10:2] ? regs__384 : _GEN_916; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_918 = 9'h181 == bpuUpdateReq_pc[10:2] ? regs__385 : _GEN_917; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_919 = 9'h182 == bpuUpdateReq_pc[10:2] ? regs__386 : _GEN_918; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_920 = 9'h183 == bpuUpdateReq_pc[10:2] ? regs__387 : _GEN_919; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_921 = 9'h184 == bpuUpdateReq_pc[10:2] ? regs__388 : _GEN_920; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_922 = 9'h185 == bpuUpdateReq_pc[10:2] ? regs__389 : _GEN_921; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_923 = 9'h186 == bpuUpdateReq_pc[10:2] ? regs__390 : _GEN_922; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_924 = 9'h187 == bpuUpdateReq_pc[10:2] ? regs__391 : _GEN_923; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_925 = 9'h188 == bpuUpdateReq_pc[10:2] ? regs__392 : _GEN_924; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_926 = 9'h189 == bpuUpdateReq_pc[10:2] ? regs__393 : _GEN_925; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_927 = 9'h18a == bpuUpdateReq_pc[10:2] ? regs__394 : _GEN_926; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_928 = 9'h18b == bpuUpdateReq_pc[10:2] ? regs__395 : _GEN_927; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_929 = 9'h18c == bpuUpdateReq_pc[10:2] ? regs__396 : _GEN_928; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_930 = 9'h18d == bpuUpdateReq_pc[10:2] ? regs__397 : _GEN_929; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_931 = 9'h18e == bpuUpdateReq_pc[10:2] ? regs__398 : _GEN_930; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_932 = 9'h18f == bpuUpdateReq_pc[10:2] ? regs__399 : _GEN_931; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_933 = 9'h190 == bpuUpdateReq_pc[10:2] ? regs__400 : _GEN_932; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_934 = 9'h191 == bpuUpdateReq_pc[10:2] ? regs__401 : _GEN_933; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_935 = 9'h192 == bpuUpdateReq_pc[10:2] ? regs__402 : _GEN_934; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_936 = 9'h193 == bpuUpdateReq_pc[10:2] ? regs__403 : _GEN_935; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_937 = 9'h194 == bpuUpdateReq_pc[10:2] ? regs__404 : _GEN_936; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_938 = 9'h195 == bpuUpdateReq_pc[10:2] ? regs__405 : _GEN_937; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_939 = 9'h196 == bpuUpdateReq_pc[10:2] ? regs__406 : _GEN_938; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_940 = 9'h197 == bpuUpdateReq_pc[10:2] ? regs__407 : _GEN_939; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_941 = 9'h198 == bpuUpdateReq_pc[10:2] ? regs__408 : _GEN_940; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_942 = 9'h199 == bpuUpdateReq_pc[10:2] ? regs__409 : _GEN_941; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_943 = 9'h19a == bpuUpdateReq_pc[10:2] ? regs__410 : _GEN_942; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_944 = 9'h19b == bpuUpdateReq_pc[10:2] ? regs__411 : _GEN_943; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_945 = 9'h19c == bpuUpdateReq_pc[10:2] ? regs__412 : _GEN_944; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_946 = 9'h19d == bpuUpdateReq_pc[10:2] ? regs__413 : _GEN_945; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_947 = 9'h19e == bpuUpdateReq_pc[10:2] ? regs__414 : _GEN_946; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_948 = 9'h19f == bpuUpdateReq_pc[10:2] ? regs__415 : _GEN_947; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_949 = 9'h1a0 == bpuUpdateReq_pc[10:2] ? regs__416 : _GEN_948; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_950 = 9'h1a1 == bpuUpdateReq_pc[10:2] ? regs__417 : _GEN_949; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_951 = 9'h1a2 == bpuUpdateReq_pc[10:2] ? regs__418 : _GEN_950; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_952 = 9'h1a3 == bpuUpdateReq_pc[10:2] ? regs__419 : _GEN_951; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_953 = 9'h1a4 == bpuUpdateReq_pc[10:2] ? regs__420 : _GEN_952; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_954 = 9'h1a5 == bpuUpdateReq_pc[10:2] ? regs__421 : _GEN_953; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_955 = 9'h1a6 == bpuUpdateReq_pc[10:2] ? regs__422 : _GEN_954; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_956 = 9'h1a7 == bpuUpdateReq_pc[10:2] ? regs__423 : _GEN_955; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_957 = 9'h1a8 == bpuUpdateReq_pc[10:2] ? regs__424 : _GEN_956; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_958 = 9'h1a9 == bpuUpdateReq_pc[10:2] ? regs__425 : _GEN_957; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_959 = 9'h1aa == bpuUpdateReq_pc[10:2] ? regs__426 : _GEN_958; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_960 = 9'h1ab == bpuUpdateReq_pc[10:2] ? regs__427 : _GEN_959; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_961 = 9'h1ac == bpuUpdateReq_pc[10:2] ? regs__428 : _GEN_960; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_962 = 9'h1ad == bpuUpdateReq_pc[10:2] ? regs__429 : _GEN_961; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_963 = 9'h1ae == bpuUpdateReq_pc[10:2] ? regs__430 : _GEN_962; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_964 = 9'h1af == bpuUpdateReq_pc[10:2] ? regs__431 : _GEN_963; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_965 = 9'h1b0 == bpuUpdateReq_pc[10:2] ? regs__432 : _GEN_964; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_966 = 9'h1b1 == bpuUpdateReq_pc[10:2] ? regs__433 : _GEN_965; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_967 = 9'h1b2 == bpuUpdateReq_pc[10:2] ? regs__434 : _GEN_966; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_968 = 9'h1b3 == bpuUpdateReq_pc[10:2] ? regs__435 : _GEN_967; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_969 = 9'h1b4 == bpuUpdateReq_pc[10:2] ? regs__436 : _GEN_968; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_970 = 9'h1b5 == bpuUpdateReq_pc[10:2] ? regs__437 : _GEN_969; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_971 = 9'h1b6 == bpuUpdateReq_pc[10:2] ? regs__438 : _GEN_970; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_972 = 9'h1b7 == bpuUpdateReq_pc[10:2] ? regs__439 : _GEN_971; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_973 = 9'h1b8 == bpuUpdateReq_pc[10:2] ? regs__440 : _GEN_972; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_974 = 9'h1b9 == bpuUpdateReq_pc[10:2] ? regs__441 : _GEN_973; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_975 = 9'h1ba == bpuUpdateReq_pc[10:2] ? regs__442 : _GEN_974; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_976 = 9'h1bb == bpuUpdateReq_pc[10:2] ? regs__443 : _GEN_975; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_977 = 9'h1bc == bpuUpdateReq_pc[10:2] ? regs__444 : _GEN_976; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_978 = 9'h1bd == bpuUpdateReq_pc[10:2] ? regs__445 : _GEN_977; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_979 = 9'h1be == bpuUpdateReq_pc[10:2] ? regs__446 : _GEN_978; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_980 = 9'h1bf == bpuUpdateReq_pc[10:2] ? regs__447 : _GEN_979; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_981 = 9'h1c0 == bpuUpdateReq_pc[10:2] ? regs__448 : _GEN_980; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_982 = 9'h1c1 == bpuUpdateReq_pc[10:2] ? regs__449 : _GEN_981; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_983 = 9'h1c2 == bpuUpdateReq_pc[10:2] ? regs__450 : _GEN_982; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_984 = 9'h1c3 == bpuUpdateReq_pc[10:2] ? regs__451 : _GEN_983; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_985 = 9'h1c4 == bpuUpdateReq_pc[10:2] ? regs__452 : _GEN_984; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_986 = 9'h1c5 == bpuUpdateReq_pc[10:2] ? regs__453 : _GEN_985; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_987 = 9'h1c6 == bpuUpdateReq_pc[10:2] ? regs__454 : _GEN_986; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_988 = 9'h1c7 == bpuUpdateReq_pc[10:2] ? regs__455 : _GEN_987; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_989 = 9'h1c8 == bpuUpdateReq_pc[10:2] ? regs__456 : _GEN_988; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_990 = 9'h1c9 == bpuUpdateReq_pc[10:2] ? regs__457 : _GEN_989; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_991 = 9'h1ca == bpuUpdateReq_pc[10:2] ? regs__458 : _GEN_990; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_992 = 9'h1cb == bpuUpdateReq_pc[10:2] ? regs__459 : _GEN_991; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_993 = 9'h1cc == bpuUpdateReq_pc[10:2] ? regs__460 : _GEN_992; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_994 = 9'h1cd == bpuUpdateReq_pc[10:2] ? regs__461 : _GEN_993; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_995 = 9'h1ce == bpuUpdateReq_pc[10:2] ? regs__462 : _GEN_994; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_996 = 9'h1cf == bpuUpdateReq_pc[10:2] ? regs__463 : _GEN_995; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_997 = 9'h1d0 == bpuUpdateReq_pc[10:2] ? regs__464 : _GEN_996; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_998 = 9'h1d1 == bpuUpdateReq_pc[10:2] ? regs__465 : _GEN_997; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_999 = 9'h1d2 == bpuUpdateReq_pc[10:2] ? regs__466 : _GEN_998; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_1000 = 9'h1d3 == bpuUpdateReq_pc[10:2] ? regs__467 : _GEN_999; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_1001 = 9'h1d4 == bpuUpdateReq_pc[10:2] ? regs__468 : _GEN_1000; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_1002 = 9'h1d5 == bpuUpdateReq_pc[10:2] ? regs__469 : _GEN_1001; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_1003 = 9'h1d6 == bpuUpdateReq_pc[10:2] ? regs__470 : _GEN_1002; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_1004 = 9'h1d7 == bpuUpdateReq_pc[10:2] ? regs__471 : _GEN_1003; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_1005 = 9'h1d8 == bpuUpdateReq_pc[10:2] ? regs__472 : _GEN_1004; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_1006 = 9'h1d9 == bpuUpdateReq_pc[10:2] ? regs__473 : _GEN_1005; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_1007 = 9'h1da == bpuUpdateReq_pc[10:2] ? regs__474 : _GEN_1006; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_1008 = 9'h1db == bpuUpdateReq_pc[10:2] ? regs__475 : _GEN_1007; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_1009 = 9'h1dc == bpuUpdateReq_pc[10:2] ? regs__476 : _GEN_1008; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_1010 = 9'h1dd == bpuUpdateReq_pc[10:2] ? regs__477 : _GEN_1009; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_1011 = 9'h1de == bpuUpdateReq_pc[10:2] ? regs__478 : _GEN_1010; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_1012 = 9'h1df == bpuUpdateReq_pc[10:2] ? regs__479 : _GEN_1011; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_1013 = 9'h1e0 == bpuUpdateReq_pc[10:2] ? regs__480 : _GEN_1012; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_1014 = 9'h1e1 == bpuUpdateReq_pc[10:2] ? regs__481 : _GEN_1013; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_1015 = 9'h1e2 == bpuUpdateReq_pc[10:2] ? regs__482 : _GEN_1014; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_1016 = 9'h1e3 == bpuUpdateReq_pc[10:2] ? regs__483 : _GEN_1015; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_1017 = 9'h1e4 == bpuUpdateReq_pc[10:2] ? regs__484 : _GEN_1016; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_1018 = 9'h1e5 == bpuUpdateReq_pc[10:2] ? regs__485 : _GEN_1017; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_1019 = 9'h1e6 == bpuUpdateReq_pc[10:2] ? regs__486 : _GEN_1018; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_1020 = 9'h1e7 == bpuUpdateReq_pc[10:2] ? regs__487 : _GEN_1019; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_1021 = 9'h1e8 == bpuUpdateReq_pc[10:2] ? regs__488 : _GEN_1020; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_1022 = 9'h1e9 == bpuUpdateReq_pc[10:2] ? regs__489 : _GEN_1021; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_1023 = 9'h1ea == bpuUpdateReq_pc[10:2] ? regs__490 : _GEN_1022; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_1024 = 9'h1eb == bpuUpdateReq_pc[10:2] ? regs__491 : _GEN_1023; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_1025 = 9'h1ec == bpuUpdateReq_pc[10:2] ? regs__492 : _GEN_1024; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_1026 = 9'h1ed == bpuUpdateReq_pc[10:2] ? regs__493 : _GEN_1025; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_1027 = 9'h1ee == bpuUpdateReq_pc[10:2] ? regs__494 : _GEN_1026; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_1028 = 9'h1ef == bpuUpdateReq_pc[10:2] ? regs__495 : _GEN_1027; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_1029 = 9'h1f0 == bpuUpdateReq_pc[10:2] ? regs__496 : _GEN_1028; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_1030 = 9'h1f1 == bpuUpdateReq_pc[10:2] ? regs__497 : _GEN_1029; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_1031 = 9'h1f2 == bpuUpdateReq_pc[10:2] ? regs__498 : _GEN_1030; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_1032 = 9'h1f3 == bpuUpdateReq_pc[10:2] ? regs__499 : _GEN_1031; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_1033 = 9'h1f4 == bpuUpdateReq_pc[10:2] ? regs__500 : _GEN_1032; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_1034 = 9'h1f5 == bpuUpdateReq_pc[10:2] ? regs__501 : _GEN_1033; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_1035 = 9'h1f6 == bpuUpdateReq_pc[10:2] ? regs__502 : _GEN_1034; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_1036 = 9'h1f7 == bpuUpdateReq_pc[10:2] ? regs__503 : _GEN_1035; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_1037 = 9'h1f8 == bpuUpdateReq_pc[10:2] ? regs__504 : _GEN_1036; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_1038 = 9'h1f9 == bpuUpdateReq_pc[10:2] ? regs__505 : _GEN_1037; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_1039 = 9'h1fa == bpuUpdateReq_pc[10:2] ? regs__506 : _GEN_1038; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  wire [1:0] _GEN_1040 = 9'h1fb == bpuUpdateReq_pc[10:2] ? regs__507 : _GEN_1039; // @[src/main/scala/nutcore/frontend/BPU.scala 389:{20,20}]
  reg  reqLatch_valid; // @[src/main/scala/nutcore/frontend/BPU.scala 390:25]
  reg [38:0] reqLatch_pc; // @[src/main/scala/nutcore/frontend/BPU.scala 390:25]
  reg  reqLatch_actualTaken; // @[src/main/scala/nutcore/frontend/BPU.scala 390:25]
  reg [6:0] reqLatch_fuOpType; // @[src/main/scala/nutcore/frontend/BPU.scala 390:25]
  wire  _T_43 = ~reqLatch_fuOpType[3]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 63:30]
  wire [1:0] _newCnt_T_1 = cnt + 2'h1; // @[src/main/scala/nutcore/frontend/BPU.scala 393:33]
  wire [1:0] _newCnt_T_3 = cnt - 2'h1; // @[src/main/scala/nutcore/frontend/BPU.scala 393:44]
  wire [1:0] newCnt = reqLatch_actualTaken ? _newCnt_T_1 : _newCnt_T_3; // @[src/main/scala/nutcore/frontend/BPU.scala 393:21]
  wire  wen = reqLatch_actualTaken & cnt != 2'h3 | ~reqLatch_actualTaken & cnt != 2'h0; // @[src/main/scala/nutcore/frontend/BPU.scala 394:44]
  wire [3:0] _T_50 = sp_value + 4'h1; // @[src/main/scala/nutcore/frontend/BPU.scala 404:26]
  wire [38:0] _T_52 = bpuUpdateReq_pc + 39'h2; // @[src/main/scala/nutcore/frontend/BPU.scala 404:55]
  wire [38:0] _T_54 = bpuUpdateReq_pc + 39'h4; // @[src/main/scala/nutcore/frontend/BPU.scala 404:69]
  wire [38:0] _T_55 = bpuUpdateReq_isRVC ? _T_52 : _T_54; // @[src/main/scala/nutcore/frontend/BPU.scala 404:36]
  wire  _T_57 = sp_value == 4'h0; // @[src/main/scala/nutcore/frontend/BPU.scala 409:21]
  wire [3:0] _value_T_4 = sp_value - 4'h1; // @[src/main/scala/nutcore/frontend/BPU.scala 412:53]
  wire [3:0] _value_T_5 = _T_57 ? 4'h0 : _value_T_4; // @[src/main/scala/nutcore/frontend/BPU.scala 412:22]
  wire [1:0] btbRead__type = btb_io_r_resp_data_0__type; // @[src/main/scala/nutcore/frontend/BPU.scala 315:21 316:11]
  wire [38:0] btbRead_target = btb_io_r_resp_data_0_target; // @[src/main/scala/nutcore/frontend/BPU.scala 315:21 316:11]
  wire [3:0] _io_brIdx_T_2 = {1'h1,crosslineJump,_T_20}; // @[src/main/scala/nutcore/frontend/BPU.scala 419:35]
  wire [3:0] _GEN_2632 = {{1'd0}, btbRead_brIdx}; // @[src/main/scala/nutcore/frontend/BPU.scala 419:30]
  wire [3:0] _io_brIdx_T_3 = _GEN_2632 & _io_brIdx_T_2; // @[src/main/scala/nutcore/frontend/BPU.scala 419:30]
  wire  _io_out_valid_T_3 = btbRead__type == 2'h0 ? phtTaken : rasTarget != 39'h0; // @[src/main/scala/nutcore/frontend/BPU.scala 420:32]
  SRAMTemplate btb ( // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
    .clock(btb_clock),
    .reset(btb_reset),
    .io_r_req_ready(btb_io_r_req_ready),
    .io_r_req_valid(btb_io_r_req_valid),
    .io_r_req_bits_setIdx(btb_io_r_req_bits_setIdx),
    .io_r_resp_data_0_tag(btb_io_r_resp_data_0_tag),
    .io_r_resp_data_0__type(btb_io_r_resp_data_0__type),
    .io_r_resp_data_0_target(btb_io_r_resp_data_0_target),
    .io_r_resp_data_0_brIdx(btb_io_r_resp_data_0_brIdx),
    .io_r_resp_data_0_valid(btb_io_r_resp_data_0_valid),
    .io_w_req_valid(btb_io_w_req_valid),
    .io_w_req_bits_setIdx(btb_io_w_req_bits_setIdx),
    .io_w_req_bits_data_tag(btb_io_w_req_bits_data_tag),
    .io_w_req_bits_data__type(btb_io_w_req_bits_data__type),
    .io_w_req_bits_data_target(btb_io_w_req_bits_data_target),
    .io_w_req_bits_data_brIdx(btb_io_w_req_bits_data_brIdx)
  );
  assign io_out_target = btbRead__type == 2'h3 ? rasTarget : btbRead_target; // @[src/main/scala/nutcore/frontend/BPU.scala 416:23]
  assign io_out_valid = btbHit & _io_out_valid_T_3; // @[src/main/scala/nutcore/frontend/BPU.scala 420:26]
  assign io_brIdx = _io_brIdx_T_3[2:0]; // @[src/main/scala/nutcore/frontend/BPU.scala 419:13]
  assign io_crosslineJump = btbRead_brIdx[2] & btbHit; // @[src/main/scala/nutcore/frontend/BPU.scala 327:40]
  assign btb_clock = clock;
  assign btb_reset = reset | (MOUFlushICache | MOUFlushTLB); // @[src/main/scala/nutcore/frontend/BPU.scala 308:29]
  assign btb_io_r_req_valid = io_in_pc_valid; // @[src/main/scala/nutcore/frontend/BPU.scala 311:22]
  assign btb_io_r_req_bits_setIdx = io_in_pc_bits[10:2]; // @[src/main/scala/nutcore/frontend/BPU.scala 35:65]
  assign btb_io_w_req_valid = bpuUpdateReq_isMissPredict & bpuUpdateReq_valid; // @[src/main/scala/nutcore/frontend/BPU.scala 375:43]
  assign btb_io_w_req_bits_setIdx = bpuUpdateReq_pc[10:2]; // @[src/main/scala/nutcore/frontend/BPU.scala 35:65]
  assign btb_io_w_req_bits_data_tag = bpuUpdateReq_pc[38:11]; // @[src/main/scala/nutcore/frontend/BPU.scala 35:65]
  assign btb_io_w_req_bits_data__type = bpuUpdateReq_btbType; // @[src/main/scala/nutcore/frontend/BPU.scala 349:21]
  assign btb_io_w_req_bits_data_target = bpuUpdateReq_actualTarget; // @[src/main/scala/nutcore/frontend/BPU.scala 349:21]
  assign btb_io_w_req_bits_data_brIdx = {btbWrite_brIdx_hi,_T_35}; // @[src/main/scala/nutcore/frontend/BPU.scala 367:24]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      flush <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      flush <= _GEN_1;
    end
    if (io_in_pc_valid) begin // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
      pcLatch <= io_in_pc_bits; // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    if (reset) begin // @[src/main/scala/nutcore/frontend/BPU.scala 320:93]
      btbHit_REG <= 1'h0; // @[src/main/scala/nutcore/frontend/BPU.scala 320:93]
    end else begin
      btbHit_REG <= _btbHit_T_7; // @[src/main/scala/nutcore/frontend/BPU.scala 320:93]
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__0 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h0 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__0 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__1 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__1 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__2 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h2 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__2 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__3 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h3 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__3 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__4 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h4 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__4 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__5 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h5 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__5 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__6 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h6 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__6 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__7 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h7 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__7 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__8 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h8 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__8 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__9 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h9 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__9 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__10 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'ha == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__10 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__11 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hb == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__11 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__12 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hc == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__12 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__13 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hd == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__13 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__14 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'he == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__14 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__15 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hf == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__15 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__16 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h10 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__16 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__17 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h11 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__17 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__18 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h12 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__18 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__19 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h13 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__19 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__20 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h14 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__20 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__21 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h15 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__21 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__22 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h16 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__22 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__23 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h17 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__23 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__24 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h18 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__24 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__25 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h19 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__25 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__26 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1a == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__26 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__27 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1b == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__27 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__28 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1c == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__28 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__29 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1d == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__29 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__30 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1e == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__30 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__31 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1f == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__31 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__32 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h20 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__32 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__33 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h21 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__33 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__34 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h22 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__34 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__35 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h23 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__35 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__36 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h24 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__36 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__37 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h25 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__37 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__38 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h26 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__38 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__39 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h27 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__39 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__40 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h28 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__40 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__41 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h29 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__41 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__42 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h2a == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__42 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__43 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h2b == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__43 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__44 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h2c == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__44 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__45 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h2d == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__45 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__46 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h2e == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__46 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__47 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h2f == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__47 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__48 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h30 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__48 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__49 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h31 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__49 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__50 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h32 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__50 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__51 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h33 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__51 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__52 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h34 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__52 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__53 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h35 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__53 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__54 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h36 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__54 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__55 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h37 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__55 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__56 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h38 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__56 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__57 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h39 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__57 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__58 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h3a == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__58 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__59 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h3b == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__59 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__60 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h3c == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__60 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__61 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h3d == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__61 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__62 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h3e == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__62 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__63 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h3f == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__63 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__64 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h40 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__64 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__65 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h41 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__65 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__66 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h42 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__66 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__67 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h43 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__67 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__68 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h44 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__68 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__69 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h45 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__69 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__70 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h46 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__70 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__71 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h47 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__71 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__72 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h48 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__72 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__73 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h49 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__73 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__74 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h4a == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__74 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__75 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h4b == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__75 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__76 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h4c == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__76 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__77 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h4d == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__77 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__78 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h4e == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__78 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__79 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h4f == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__79 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__80 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h50 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__80 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__81 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h51 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__81 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__82 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h52 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__82 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__83 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h53 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__83 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__84 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h54 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__84 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__85 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h55 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__85 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__86 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h56 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__86 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__87 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h57 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__87 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__88 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h58 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__88 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__89 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h59 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__89 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__90 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h5a == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__90 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__91 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h5b == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__91 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__92 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h5c == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__92 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__93 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h5d == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__93 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__94 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h5e == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__94 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__95 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h5f == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__95 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__96 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h60 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__96 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__97 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h61 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__97 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__98 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h62 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__98 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__99 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h63 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__99 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__100 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h64 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__100 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__101 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h65 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__101 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__102 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h66 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__102 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__103 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h67 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__103 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__104 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h68 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__104 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__105 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h69 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__105 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__106 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h6a == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__106 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__107 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h6b == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__107 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__108 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h6c == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__108 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__109 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h6d == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__109 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__110 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h6e == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__110 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__111 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h6f == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__111 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__112 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h70 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__112 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__113 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h71 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__113 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__114 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h72 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__114 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__115 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h73 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__115 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__116 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h74 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__116 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__117 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h75 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__117 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__118 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h76 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__118 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__119 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h77 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__119 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__120 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h78 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__120 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__121 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h79 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__121 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__122 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h7a == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__122 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__123 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h7b == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__123 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__124 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h7c == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__124 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__125 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h7d == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__125 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__126 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h7e == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__126 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__127 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h7f == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__127 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__128 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h80 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__128 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__129 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h81 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__129 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__130 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h82 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__130 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__131 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h83 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__131 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__132 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h84 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__132 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__133 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h85 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__133 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__134 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h86 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__134 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__135 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h87 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__135 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__136 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h88 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__136 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__137 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h89 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__137 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__138 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h8a == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__138 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__139 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h8b == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__139 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__140 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h8c == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__140 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__141 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h8d == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__141 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__142 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h8e == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__142 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__143 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h8f == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__143 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__144 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h90 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__144 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__145 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h91 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__145 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__146 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h92 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__146 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__147 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h93 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__147 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__148 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h94 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__148 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__149 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h95 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__149 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__150 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h96 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__150 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__151 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h97 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__151 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__152 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h98 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__152 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__153 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h99 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__153 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__154 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h9a == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__154 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__155 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h9b == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__155 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__156 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h9c == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__156 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__157 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h9d == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__157 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__158 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h9e == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__158 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__159 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h9f == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__159 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__160 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'ha0 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__160 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__161 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'ha1 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__161 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__162 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'ha2 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__162 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__163 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'ha3 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__163 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__164 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'ha4 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__164 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__165 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'ha5 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__165 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__166 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'ha6 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__166 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__167 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'ha7 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__167 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__168 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'ha8 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__168 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__169 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'ha9 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__169 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__170 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'haa == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__170 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__171 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hab == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__171 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__172 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hac == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__172 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__173 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'had == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__173 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__174 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hae == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__174 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__175 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'haf == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__175 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__176 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hb0 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__176 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__177 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hb1 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__177 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__178 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hb2 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__178 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__179 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hb3 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__179 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__180 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hb4 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__180 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__181 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hb5 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__181 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__182 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hb6 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__182 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__183 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hb7 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__183 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__184 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hb8 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__184 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__185 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hb9 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__185 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__186 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hba == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__186 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__187 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hbb == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__187 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__188 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hbc == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__188 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__189 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hbd == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__189 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__190 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hbe == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__190 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__191 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hbf == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__191 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__192 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hc0 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__192 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__193 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hc1 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__193 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__194 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hc2 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__194 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__195 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hc3 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__195 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__196 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hc4 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__196 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__197 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hc5 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__197 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__198 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hc6 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__198 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__199 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hc7 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__199 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__200 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hc8 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__200 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__201 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hc9 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__201 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__202 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hca == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__202 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__203 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hcb == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__203 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__204 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hcc == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__204 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__205 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hcd == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__205 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__206 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hce == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__206 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__207 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hcf == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__207 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__208 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hd0 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__208 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__209 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hd1 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__209 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__210 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hd2 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__210 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__211 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hd3 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__211 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__212 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hd4 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__212 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__213 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hd5 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__213 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__214 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hd6 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__214 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__215 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hd7 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__215 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__216 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hd8 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__216 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__217 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hd9 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__217 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__218 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hda == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__218 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__219 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hdb == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__219 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__220 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hdc == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__220 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__221 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hdd == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__221 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__222 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hde == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__222 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__223 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hdf == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__223 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__224 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'he0 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__224 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__225 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'he1 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__225 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__226 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'he2 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__226 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__227 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'he3 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__227 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__228 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'he4 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__228 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__229 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'he5 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__229 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__230 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'he6 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__230 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__231 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'he7 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__231 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__232 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'he8 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__232 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__233 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'he9 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__233 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__234 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hea == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__234 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__235 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'heb == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__235 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__236 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hec == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__236 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__237 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hed == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__237 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__238 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hee == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__238 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__239 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hef == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__239 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__240 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hf0 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__240 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__241 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hf1 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__241 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__242 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hf2 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__242 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__243 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hf3 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__243 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__244 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hf4 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__244 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__245 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hf5 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__245 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__246 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hf6 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__246 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__247 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hf7 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__247 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__248 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hf8 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__248 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__249 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hf9 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__249 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__250 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hfa == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__250 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__251 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hfb == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__251 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__252 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hfc == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__252 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__253 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hfd == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__253 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__254 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hfe == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__254 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__255 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'hff == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__255 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__256 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h100 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__256 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__257 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h101 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__257 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__258 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h102 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__258 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__259 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h103 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__259 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__260 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h104 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__260 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__261 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h105 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__261 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__262 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h106 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__262 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__263 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h107 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__263 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__264 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h108 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__264 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__265 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h109 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__265 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__266 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h10a == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__266 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__267 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h10b == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__267 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__268 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h10c == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__268 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__269 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h10d == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__269 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__270 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h10e == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__270 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__271 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h10f == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__271 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__272 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h110 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__272 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__273 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h111 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__273 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__274 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h112 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__274 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__275 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h113 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__275 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__276 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h114 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__276 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__277 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h115 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__277 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__278 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h116 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__278 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__279 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h117 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__279 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__280 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h118 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__280 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__281 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h119 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__281 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__282 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h11a == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__282 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__283 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h11b == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__283 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__284 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h11c == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__284 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__285 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h11d == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__285 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__286 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h11e == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__286 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__287 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h11f == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__287 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__288 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h120 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__288 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__289 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h121 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__289 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__290 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h122 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__290 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__291 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h123 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__291 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__292 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h124 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__292 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__293 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h125 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__293 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__294 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h126 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__294 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__295 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h127 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__295 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__296 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h128 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__296 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__297 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h129 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__297 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__298 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h12a == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__298 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__299 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h12b == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__299 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__300 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h12c == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__300 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__301 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h12d == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__301 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__302 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h12e == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__302 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__303 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h12f == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__303 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__304 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h130 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__304 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__305 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h131 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__305 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__306 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h132 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__306 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__307 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h133 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__307 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__308 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h134 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__308 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__309 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h135 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__309 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__310 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h136 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__310 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__311 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h137 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__311 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__312 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h138 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__312 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__313 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h139 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__313 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__314 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h13a == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__314 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__315 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h13b == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__315 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__316 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h13c == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__316 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__317 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h13d == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__317 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__318 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h13e == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__318 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__319 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h13f == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__319 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__320 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h140 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__320 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__321 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h141 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__321 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__322 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h142 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__322 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__323 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h143 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__323 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__324 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h144 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__324 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__325 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h145 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__325 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__326 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h146 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__326 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__327 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h147 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__327 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__328 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h148 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__328 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__329 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h149 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__329 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__330 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h14a == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__330 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__331 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h14b == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__331 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__332 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h14c == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__332 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__333 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h14d == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__333 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__334 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h14e == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__334 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__335 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h14f == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__335 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__336 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h150 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__336 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__337 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h151 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__337 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__338 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h152 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__338 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__339 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h153 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__339 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__340 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h154 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__340 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__341 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h155 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__341 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__342 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h156 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__342 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__343 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h157 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__343 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__344 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h158 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__344 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__345 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h159 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__345 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__346 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h15a == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__346 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__347 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h15b == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__347 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__348 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h15c == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__348 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__349 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h15d == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__349 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__350 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h15e == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__350 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__351 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h15f == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__351 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__352 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h160 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__352 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__353 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h161 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__353 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__354 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h162 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__354 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__355 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h163 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__355 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__356 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h164 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__356 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__357 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h165 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__357 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__358 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h166 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__358 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__359 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h167 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__359 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__360 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h168 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__360 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__361 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h169 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__361 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__362 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h16a == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__362 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__363 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h16b == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__363 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__364 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h16c == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__364 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__365 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h16d == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__365 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__366 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h16e == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__366 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__367 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h16f == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__367 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__368 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h170 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__368 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__369 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h171 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__369 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__370 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h172 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__370 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__371 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h173 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__371 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__372 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h174 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__372 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__373 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h175 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__373 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__374 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h176 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__374 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__375 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h177 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__375 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__376 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h178 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__376 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__377 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h179 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__377 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__378 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h17a == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__378 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__379 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h17b == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__379 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__380 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h17c == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__380 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__381 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h17d == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__381 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__382 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h17e == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__382 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__383 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h17f == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__383 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__384 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h180 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__384 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__385 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h181 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__385 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__386 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h182 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__386 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__387 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h183 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__387 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__388 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h184 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__388 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__389 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h185 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__389 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__390 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h186 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__390 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__391 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h187 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__391 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__392 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h188 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__392 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__393 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h189 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__393 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__394 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h18a == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__394 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__395 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h18b == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__395 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__396 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h18c == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__396 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__397 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h18d == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__397 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__398 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h18e == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__398 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__399 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h18f == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__399 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__400 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h190 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__400 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__401 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h191 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__401 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__402 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h192 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__402 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__403 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h193 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__403 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__404 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h194 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__404 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__405 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h195 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__405 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__406 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h196 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__406 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__407 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h197 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__407 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__408 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h198 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__408 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__409 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h199 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__409 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__410 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h19a == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__410 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__411 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h19b == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__411 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__412 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h19c == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__412 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__413 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h19d == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__413 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__414 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h19e == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__414 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__415 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h19f == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__415 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__416 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1a0 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__416 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__417 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1a1 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__417 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__418 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1a2 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__418 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__419 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1a3 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__419 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__420 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1a4 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__420 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__421 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1a5 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__421 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__422 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1a6 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__422 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__423 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1a7 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__423 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__424 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1a8 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__424 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__425 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1a9 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__425 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__426 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1aa == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__426 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__427 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1ab == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__427 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__428 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1ac == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__428 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__429 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1ad == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__429 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__430 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1ae == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__430 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__431 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1af == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__431 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__432 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1b0 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__432 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__433 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1b1 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__433 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__434 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1b2 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__434 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__435 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1b3 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__435 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__436 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1b4 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__436 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__437 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1b5 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__437 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__438 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1b6 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__438 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__439 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1b7 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__439 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__440 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1b8 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__440 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__441 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1b9 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__441 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__442 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1ba == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__442 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__443 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1bb == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__443 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__444 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1bc == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__444 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__445 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1bd == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__445 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__446 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1be == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__446 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__447 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1bf == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__447 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__448 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1c0 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__448 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__449 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1c1 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__449 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__450 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1c2 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__450 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__451 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1c3 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__451 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__452 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1c4 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__452 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__453 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1c5 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__453 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__454 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1c6 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__454 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__455 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1c7 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__455 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__456 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1c8 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__456 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__457 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1c9 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__457 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__458 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1ca == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__458 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__459 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1cb == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__459 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__460 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1cc == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__460 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__461 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1cd == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__461 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__462 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1ce == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__462 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__463 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1cf == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__463 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__464 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1d0 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__464 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__465 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1d1 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__465 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__466 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1d2 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__466 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__467 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1d3 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__467 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__468 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1d4 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__468 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__469 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1d5 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__469 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__470 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1d6 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__470 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__471 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1d7 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__471 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__472 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1d8 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__472 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__473 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1d9 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__473 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__474 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1da == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__474 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__475 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1db == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__475 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__476 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1dc == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__476 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__477 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1dd == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__477 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__478 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1de == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__478 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__479 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1df == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__479 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__480 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1e0 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__480 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__481 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1e1 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__481 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__482 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1e2 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__482 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__483 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1e3 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__483 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__484 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1e4 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__484 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__485 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1e5 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__485 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__486 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1e6 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__486 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__487 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1e7 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__487 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__488 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1e8 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__488 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__489 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1e9 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__489 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__490 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1ea == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__490 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__491 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1eb == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__491 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__492 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1ec == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__492 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__493 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1ed == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__493 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__494 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1ee == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__494 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__495 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1ef == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__495 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__496 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1f0 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__496 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__497 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1f1 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__497 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__498 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1f2 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__498 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__499 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1f3 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__499 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__500 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1f4 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__500 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__501 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1f5 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__501 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__502 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1f6 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__502 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__503 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1f7 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__503 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__504 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1f8 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__504 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__505 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1f9 == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__505 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__506 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1fa == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__506 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__507 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1fb == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__507 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__508 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1fc == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__508 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__509 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1fd == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__509 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__510 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1fe == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__510 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs__511 <= 2'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (reqLatch_valid & _T_43) begin // @[src/main/scala/nutcore/frontend/BPU.scala 391:66]
      if (wen) begin // @[src/main/scala/nutcore/frontend/BPU.scala 395:16]
        if (9'h1ff == reqLatch_pc[10:2]) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs__511 <= newCnt; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (io_in_pc_valid) begin // @[src/main/scala/nutcore/frontend/BPU.scala 337:27]
      phtTaken <= _GEN_514[1]; // @[src/main/scala/nutcore/frontend/BPU.scala 337:27]
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_1_0 <= 39'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (bpuUpdateReq_valid) begin // @[src/main/scala/nutcore/frontend/BPU.scala 402:20]
      if (bpuUpdateReq_fuOpType == 7'h5c) begin // @[src/main/scala/nutcore/frontend/BPU.scala 403:45]
        if (4'h0 == _T_50) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs_1_0 <= _T_55; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_1_1 <= 39'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (bpuUpdateReq_valid) begin // @[src/main/scala/nutcore/frontend/BPU.scala 402:20]
      if (bpuUpdateReq_fuOpType == 7'h5c) begin // @[src/main/scala/nutcore/frontend/BPU.scala 403:45]
        if (4'h1 == _T_50) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs_1_1 <= _T_55; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_1_2 <= 39'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (bpuUpdateReq_valid) begin // @[src/main/scala/nutcore/frontend/BPU.scala 402:20]
      if (bpuUpdateReq_fuOpType == 7'h5c) begin // @[src/main/scala/nutcore/frontend/BPU.scala 403:45]
        if (4'h2 == _T_50) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs_1_2 <= _T_55; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_1_3 <= 39'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (bpuUpdateReq_valid) begin // @[src/main/scala/nutcore/frontend/BPU.scala 402:20]
      if (bpuUpdateReq_fuOpType == 7'h5c) begin // @[src/main/scala/nutcore/frontend/BPU.scala 403:45]
        if (4'h3 == _T_50) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs_1_3 <= _T_55; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_1_4 <= 39'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (bpuUpdateReq_valid) begin // @[src/main/scala/nutcore/frontend/BPU.scala 402:20]
      if (bpuUpdateReq_fuOpType == 7'h5c) begin // @[src/main/scala/nutcore/frontend/BPU.scala 403:45]
        if (4'h4 == _T_50) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs_1_4 <= _T_55; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_1_5 <= 39'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (bpuUpdateReq_valid) begin // @[src/main/scala/nutcore/frontend/BPU.scala 402:20]
      if (bpuUpdateReq_fuOpType == 7'h5c) begin // @[src/main/scala/nutcore/frontend/BPU.scala 403:45]
        if (4'h5 == _T_50) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs_1_5 <= _T_55; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_1_6 <= 39'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (bpuUpdateReq_valid) begin // @[src/main/scala/nutcore/frontend/BPU.scala 402:20]
      if (bpuUpdateReq_fuOpType == 7'h5c) begin // @[src/main/scala/nutcore/frontend/BPU.scala 403:45]
        if (4'h6 == _T_50) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs_1_6 <= _T_55; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_1_7 <= 39'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (bpuUpdateReq_valid) begin // @[src/main/scala/nutcore/frontend/BPU.scala 402:20]
      if (bpuUpdateReq_fuOpType == 7'h5c) begin // @[src/main/scala/nutcore/frontend/BPU.scala 403:45]
        if (4'h7 == _T_50) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs_1_7 <= _T_55; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_1_8 <= 39'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (bpuUpdateReq_valid) begin // @[src/main/scala/nutcore/frontend/BPU.scala 402:20]
      if (bpuUpdateReq_fuOpType == 7'h5c) begin // @[src/main/scala/nutcore/frontend/BPU.scala 403:45]
        if (4'h8 == _T_50) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs_1_8 <= _T_55; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_1_9 <= 39'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (bpuUpdateReq_valid) begin // @[src/main/scala/nutcore/frontend/BPU.scala 402:20]
      if (bpuUpdateReq_fuOpType == 7'h5c) begin // @[src/main/scala/nutcore/frontend/BPU.scala 403:45]
        if (4'h9 == _T_50) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs_1_9 <= _T_55; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_1_10 <= 39'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (bpuUpdateReq_valid) begin // @[src/main/scala/nutcore/frontend/BPU.scala 402:20]
      if (bpuUpdateReq_fuOpType == 7'h5c) begin // @[src/main/scala/nutcore/frontend/BPU.scala 403:45]
        if (4'ha == _T_50) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs_1_10 <= _T_55; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_1_11 <= 39'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (bpuUpdateReq_valid) begin // @[src/main/scala/nutcore/frontend/BPU.scala 402:20]
      if (bpuUpdateReq_fuOpType == 7'h5c) begin // @[src/main/scala/nutcore/frontend/BPU.scala 403:45]
        if (4'hb == _T_50) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs_1_11 <= _T_55; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_1_12 <= 39'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (bpuUpdateReq_valid) begin // @[src/main/scala/nutcore/frontend/BPU.scala 402:20]
      if (bpuUpdateReq_fuOpType == 7'h5c) begin // @[src/main/scala/nutcore/frontend/BPU.scala 403:45]
        if (4'hc == _T_50) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs_1_12 <= _T_55; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_1_13 <= 39'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (bpuUpdateReq_valid) begin // @[src/main/scala/nutcore/frontend/BPU.scala 402:20]
      if (bpuUpdateReq_fuOpType == 7'h5c) begin // @[src/main/scala/nutcore/frontend/BPU.scala 403:45]
        if (4'hd == _T_50) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs_1_13 <= _T_55; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_1_14 <= 39'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (bpuUpdateReq_valid) begin // @[src/main/scala/nutcore/frontend/BPU.scala 402:20]
      if (bpuUpdateReq_fuOpType == 7'h5c) begin // @[src/main/scala/nutcore/frontend/BPU.scala 403:45]
        if (4'he == _T_50) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs_1_14 <= _T_55; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_1_15 <= 39'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (bpuUpdateReq_valid) begin // @[src/main/scala/nutcore/frontend/BPU.scala 402:20]
      if (bpuUpdateReq_fuOpType == 7'h5c) begin // @[src/main/scala/nutcore/frontend/BPU.scala 403:45]
        if (4'hf == _T_50) begin // @[src/main/scala/utils/RegMem.scala 13:15]
          regs_1_15 <= _T_55; // @[src/main/scala/utils/RegMem.scala 13:15]
        end
      end
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      sp_value <= 4'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (bpuUpdateReq_valid) begin // @[src/main/scala/nutcore/frontend/BPU.scala 402:20]
      if (bpuUpdateReq_fuOpType == 7'h5c) begin // @[src/main/scala/nutcore/frontend/BPU.scala 403:45]
        sp_value <= _T_50; // @[src/main/scala/nutcore/frontend/BPU.scala 406:16]
      end else if (bpuUpdateReq_fuOpType == 7'h5e) begin // @[src/main/scala/nutcore/frontend/BPU.scala 408:48]
        sp_value <= _value_T_5; // @[src/main/scala/nutcore/frontend/BPU.scala 412:16]
      end
    end
    if (io_in_pc_valid) begin // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
      if (4'hf == sp_value) begin // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
        rasTarget <= regs_1_15; // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
      end else if (4'he == sp_value) begin // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
        rasTarget <= regs_1_14; // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
      end else if (4'hd == sp_value) begin // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
        rasTarget <= regs_1_13; // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
      end else begin
        rasTarget <= _GEN_528;
      end
    end
    if (9'h1ff == bpuUpdateReq_pc[10:2]) begin // @[src/main/scala/nutcore/frontend/BPU.scala 389:20]
      cnt <= regs__511; // @[src/main/scala/nutcore/frontend/BPU.scala 389:20]
    end else if (9'h1fe == bpuUpdateReq_pc[10:2]) begin // @[src/main/scala/nutcore/frontend/BPU.scala 389:20]
      cnt <= regs__510; // @[src/main/scala/nutcore/frontend/BPU.scala 389:20]
    end else if (9'h1fd == bpuUpdateReq_pc[10:2]) begin // @[src/main/scala/nutcore/frontend/BPU.scala 389:20]
      cnt <= regs__509; // @[src/main/scala/nutcore/frontend/BPU.scala 389:20]
    end else if (9'h1fc == bpuUpdateReq_pc[10:2]) begin // @[src/main/scala/nutcore/frontend/BPU.scala 389:20]
      cnt <= regs__508; // @[src/main/scala/nutcore/frontend/BPU.scala 389:20]
    end else begin
      cnt <= _GEN_1040;
    end
    reqLatch_valid <= bpuUpdateReq_valid; // @[src/main/scala/nutcore/frontend/BPU.scala 349:21]
    reqLatch_pc <= bpuUpdateReq_pc; // @[src/main/scala/nutcore/frontend/BPU.scala 349:21]
    reqLatch_actualTaken <= bpuUpdateReq_actualTaken; // @[src/main/scala/nutcore/frontend/BPU.scala 349:21]
    reqLatch_fuOpType <= bpuUpdateReq_fuOpType; // @[src/main/scala/nutcore/frontend/BPU.scala 349:21]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  flush = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  pcLatch = _RAND_1[38:0];
  _RAND_2 = {1{`RANDOM}};
  btbHit_REG = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  regs__0 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  regs__1 = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  regs__2 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  regs__3 = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  regs__4 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  regs__5 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  regs__6 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  regs__7 = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  regs__8 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  regs__9 = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  regs__10 = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  regs__11 = _RAND_14[1:0];
  _RAND_15 = {1{`RANDOM}};
  regs__12 = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  regs__13 = _RAND_16[1:0];
  _RAND_17 = {1{`RANDOM}};
  regs__14 = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  regs__15 = _RAND_18[1:0];
  _RAND_19 = {1{`RANDOM}};
  regs__16 = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  regs__17 = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  regs__18 = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  regs__19 = _RAND_22[1:0];
  _RAND_23 = {1{`RANDOM}};
  regs__20 = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  regs__21 = _RAND_24[1:0];
  _RAND_25 = {1{`RANDOM}};
  regs__22 = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  regs__23 = _RAND_26[1:0];
  _RAND_27 = {1{`RANDOM}};
  regs__24 = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  regs__25 = _RAND_28[1:0];
  _RAND_29 = {1{`RANDOM}};
  regs__26 = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  regs__27 = _RAND_30[1:0];
  _RAND_31 = {1{`RANDOM}};
  regs__28 = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  regs__29 = _RAND_32[1:0];
  _RAND_33 = {1{`RANDOM}};
  regs__30 = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  regs__31 = _RAND_34[1:0];
  _RAND_35 = {1{`RANDOM}};
  regs__32 = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  regs__33 = _RAND_36[1:0];
  _RAND_37 = {1{`RANDOM}};
  regs__34 = _RAND_37[1:0];
  _RAND_38 = {1{`RANDOM}};
  regs__35 = _RAND_38[1:0];
  _RAND_39 = {1{`RANDOM}};
  regs__36 = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  regs__37 = _RAND_40[1:0];
  _RAND_41 = {1{`RANDOM}};
  regs__38 = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  regs__39 = _RAND_42[1:0];
  _RAND_43 = {1{`RANDOM}};
  regs__40 = _RAND_43[1:0];
  _RAND_44 = {1{`RANDOM}};
  regs__41 = _RAND_44[1:0];
  _RAND_45 = {1{`RANDOM}};
  regs__42 = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  regs__43 = _RAND_46[1:0];
  _RAND_47 = {1{`RANDOM}};
  regs__44 = _RAND_47[1:0];
  _RAND_48 = {1{`RANDOM}};
  regs__45 = _RAND_48[1:0];
  _RAND_49 = {1{`RANDOM}};
  regs__46 = _RAND_49[1:0];
  _RAND_50 = {1{`RANDOM}};
  regs__47 = _RAND_50[1:0];
  _RAND_51 = {1{`RANDOM}};
  regs__48 = _RAND_51[1:0];
  _RAND_52 = {1{`RANDOM}};
  regs__49 = _RAND_52[1:0];
  _RAND_53 = {1{`RANDOM}};
  regs__50 = _RAND_53[1:0];
  _RAND_54 = {1{`RANDOM}};
  regs__51 = _RAND_54[1:0];
  _RAND_55 = {1{`RANDOM}};
  regs__52 = _RAND_55[1:0];
  _RAND_56 = {1{`RANDOM}};
  regs__53 = _RAND_56[1:0];
  _RAND_57 = {1{`RANDOM}};
  regs__54 = _RAND_57[1:0];
  _RAND_58 = {1{`RANDOM}};
  regs__55 = _RAND_58[1:0];
  _RAND_59 = {1{`RANDOM}};
  regs__56 = _RAND_59[1:0];
  _RAND_60 = {1{`RANDOM}};
  regs__57 = _RAND_60[1:0];
  _RAND_61 = {1{`RANDOM}};
  regs__58 = _RAND_61[1:0];
  _RAND_62 = {1{`RANDOM}};
  regs__59 = _RAND_62[1:0];
  _RAND_63 = {1{`RANDOM}};
  regs__60 = _RAND_63[1:0];
  _RAND_64 = {1{`RANDOM}};
  regs__61 = _RAND_64[1:0];
  _RAND_65 = {1{`RANDOM}};
  regs__62 = _RAND_65[1:0];
  _RAND_66 = {1{`RANDOM}};
  regs__63 = _RAND_66[1:0];
  _RAND_67 = {1{`RANDOM}};
  regs__64 = _RAND_67[1:0];
  _RAND_68 = {1{`RANDOM}};
  regs__65 = _RAND_68[1:0];
  _RAND_69 = {1{`RANDOM}};
  regs__66 = _RAND_69[1:0];
  _RAND_70 = {1{`RANDOM}};
  regs__67 = _RAND_70[1:0];
  _RAND_71 = {1{`RANDOM}};
  regs__68 = _RAND_71[1:0];
  _RAND_72 = {1{`RANDOM}};
  regs__69 = _RAND_72[1:0];
  _RAND_73 = {1{`RANDOM}};
  regs__70 = _RAND_73[1:0];
  _RAND_74 = {1{`RANDOM}};
  regs__71 = _RAND_74[1:0];
  _RAND_75 = {1{`RANDOM}};
  regs__72 = _RAND_75[1:0];
  _RAND_76 = {1{`RANDOM}};
  regs__73 = _RAND_76[1:0];
  _RAND_77 = {1{`RANDOM}};
  regs__74 = _RAND_77[1:0];
  _RAND_78 = {1{`RANDOM}};
  regs__75 = _RAND_78[1:0];
  _RAND_79 = {1{`RANDOM}};
  regs__76 = _RAND_79[1:0];
  _RAND_80 = {1{`RANDOM}};
  regs__77 = _RAND_80[1:0];
  _RAND_81 = {1{`RANDOM}};
  regs__78 = _RAND_81[1:0];
  _RAND_82 = {1{`RANDOM}};
  regs__79 = _RAND_82[1:0];
  _RAND_83 = {1{`RANDOM}};
  regs__80 = _RAND_83[1:0];
  _RAND_84 = {1{`RANDOM}};
  regs__81 = _RAND_84[1:0];
  _RAND_85 = {1{`RANDOM}};
  regs__82 = _RAND_85[1:0];
  _RAND_86 = {1{`RANDOM}};
  regs__83 = _RAND_86[1:0];
  _RAND_87 = {1{`RANDOM}};
  regs__84 = _RAND_87[1:0];
  _RAND_88 = {1{`RANDOM}};
  regs__85 = _RAND_88[1:0];
  _RAND_89 = {1{`RANDOM}};
  regs__86 = _RAND_89[1:0];
  _RAND_90 = {1{`RANDOM}};
  regs__87 = _RAND_90[1:0];
  _RAND_91 = {1{`RANDOM}};
  regs__88 = _RAND_91[1:0];
  _RAND_92 = {1{`RANDOM}};
  regs__89 = _RAND_92[1:0];
  _RAND_93 = {1{`RANDOM}};
  regs__90 = _RAND_93[1:0];
  _RAND_94 = {1{`RANDOM}};
  regs__91 = _RAND_94[1:0];
  _RAND_95 = {1{`RANDOM}};
  regs__92 = _RAND_95[1:0];
  _RAND_96 = {1{`RANDOM}};
  regs__93 = _RAND_96[1:0];
  _RAND_97 = {1{`RANDOM}};
  regs__94 = _RAND_97[1:0];
  _RAND_98 = {1{`RANDOM}};
  regs__95 = _RAND_98[1:0];
  _RAND_99 = {1{`RANDOM}};
  regs__96 = _RAND_99[1:0];
  _RAND_100 = {1{`RANDOM}};
  regs__97 = _RAND_100[1:0];
  _RAND_101 = {1{`RANDOM}};
  regs__98 = _RAND_101[1:0];
  _RAND_102 = {1{`RANDOM}};
  regs__99 = _RAND_102[1:0];
  _RAND_103 = {1{`RANDOM}};
  regs__100 = _RAND_103[1:0];
  _RAND_104 = {1{`RANDOM}};
  regs__101 = _RAND_104[1:0];
  _RAND_105 = {1{`RANDOM}};
  regs__102 = _RAND_105[1:0];
  _RAND_106 = {1{`RANDOM}};
  regs__103 = _RAND_106[1:0];
  _RAND_107 = {1{`RANDOM}};
  regs__104 = _RAND_107[1:0];
  _RAND_108 = {1{`RANDOM}};
  regs__105 = _RAND_108[1:0];
  _RAND_109 = {1{`RANDOM}};
  regs__106 = _RAND_109[1:0];
  _RAND_110 = {1{`RANDOM}};
  regs__107 = _RAND_110[1:0];
  _RAND_111 = {1{`RANDOM}};
  regs__108 = _RAND_111[1:0];
  _RAND_112 = {1{`RANDOM}};
  regs__109 = _RAND_112[1:0];
  _RAND_113 = {1{`RANDOM}};
  regs__110 = _RAND_113[1:0];
  _RAND_114 = {1{`RANDOM}};
  regs__111 = _RAND_114[1:0];
  _RAND_115 = {1{`RANDOM}};
  regs__112 = _RAND_115[1:0];
  _RAND_116 = {1{`RANDOM}};
  regs__113 = _RAND_116[1:0];
  _RAND_117 = {1{`RANDOM}};
  regs__114 = _RAND_117[1:0];
  _RAND_118 = {1{`RANDOM}};
  regs__115 = _RAND_118[1:0];
  _RAND_119 = {1{`RANDOM}};
  regs__116 = _RAND_119[1:0];
  _RAND_120 = {1{`RANDOM}};
  regs__117 = _RAND_120[1:0];
  _RAND_121 = {1{`RANDOM}};
  regs__118 = _RAND_121[1:0];
  _RAND_122 = {1{`RANDOM}};
  regs__119 = _RAND_122[1:0];
  _RAND_123 = {1{`RANDOM}};
  regs__120 = _RAND_123[1:0];
  _RAND_124 = {1{`RANDOM}};
  regs__121 = _RAND_124[1:0];
  _RAND_125 = {1{`RANDOM}};
  regs__122 = _RAND_125[1:0];
  _RAND_126 = {1{`RANDOM}};
  regs__123 = _RAND_126[1:0];
  _RAND_127 = {1{`RANDOM}};
  regs__124 = _RAND_127[1:0];
  _RAND_128 = {1{`RANDOM}};
  regs__125 = _RAND_128[1:0];
  _RAND_129 = {1{`RANDOM}};
  regs__126 = _RAND_129[1:0];
  _RAND_130 = {1{`RANDOM}};
  regs__127 = _RAND_130[1:0];
  _RAND_131 = {1{`RANDOM}};
  regs__128 = _RAND_131[1:0];
  _RAND_132 = {1{`RANDOM}};
  regs__129 = _RAND_132[1:0];
  _RAND_133 = {1{`RANDOM}};
  regs__130 = _RAND_133[1:0];
  _RAND_134 = {1{`RANDOM}};
  regs__131 = _RAND_134[1:0];
  _RAND_135 = {1{`RANDOM}};
  regs__132 = _RAND_135[1:0];
  _RAND_136 = {1{`RANDOM}};
  regs__133 = _RAND_136[1:0];
  _RAND_137 = {1{`RANDOM}};
  regs__134 = _RAND_137[1:0];
  _RAND_138 = {1{`RANDOM}};
  regs__135 = _RAND_138[1:0];
  _RAND_139 = {1{`RANDOM}};
  regs__136 = _RAND_139[1:0];
  _RAND_140 = {1{`RANDOM}};
  regs__137 = _RAND_140[1:0];
  _RAND_141 = {1{`RANDOM}};
  regs__138 = _RAND_141[1:0];
  _RAND_142 = {1{`RANDOM}};
  regs__139 = _RAND_142[1:0];
  _RAND_143 = {1{`RANDOM}};
  regs__140 = _RAND_143[1:0];
  _RAND_144 = {1{`RANDOM}};
  regs__141 = _RAND_144[1:0];
  _RAND_145 = {1{`RANDOM}};
  regs__142 = _RAND_145[1:0];
  _RAND_146 = {1{`RANDOM}};
  regs__143 = _RAND_146[1:0];
  _RAND_147 = {1{`RANDOM}};
  regs__144 = _RAND_147[1:0];
  _RAND_148 = {1{`RANDOM}};
  regs__145 = _RAND_148[1:0];
  _RAND_149 = {1{`RANDOM}};
  regs__146 = _RAND_149[1:0];
  _RAND_150 = {1{`RANDOM}};
  regs__147 = _RAND_150[1:0];
  _RAND_151 = {1{`RANDOM}};
  regs__148 = _RAND_151[1:0];
  _RAND_152 = {1{`RANDOM}};
  regs__149 = _RAND_152[1:0];
  _RAND_153 = {1{`RANDOM}};
  regs__150 = _RAND_153[1:0];
  _RAND_154 = {1{`RANDOM}};
  regs__151 = _RAND_154[1:0];
  _RAND_155 = {1{`RANDOM}};
  regs__152 = _RAND_155[1:0];
  _RAND_156 = {1{`RANDOM}};
  regs__153 = _RAND_156[1:0];
  _RAND_157 = {1{`RANDOM}};
  regs__154 = _RAND_157[1:0];
  _RAND_158 = {1{`RANDOM}};
  regs__155 = _RAND_158[1:0];
  _RAND_159 = {1{`RANDOM}};
  regs__156 = _RAND_159[1:0];
  _RAND_160 = {1{`RANDOM}};
  regs__157 = _RAND_160[1:0];
  _RAND_161 = {1{`RANDOM}};
  regs__158 = _RAND_161[1:0];
  _RAND_162 = {1{`RANDOM}};
  regs__159 = _RAND_162[1:0];
  _RAND_163 = {1{`RANDOM}};
  regs__160 = _RAND_163[1:0];
  _RAND_164 = {1{`RANDOM}};
  regs__161 = _RAND_164[1:0];
  _RAND_165 = {1{`RANDOM}};
  regs__162 = _RAND_165[1:0];
  _RAND_166 = {1{`RANDOM}};
  regs__163 = _RAND_166[1:0];
  _RAND_167 = {1{`RANDOM}};
  regs__164 = _RAND_167[1:0];
  _RAND_168 = {1{`RANDOM}};
  regs__165 = _RAND_168[1:0];
  _RAND_169 = {1{`RANDOM}};
  regs__166 = _RAND_169[1:0];
  _RAND_170 = {1{`RANDOM}};
  regs__167 = _RAND_170[1:0];
  _RAND_171 = {1{`RANDOM}};
  regs__168 = _RAND_171[1:0];
  _RAND_172 = {1{`RANDOM}};
  regs__169 = _RAND_172[1:0];
  _RAND_173 = {1{`RANDOM}};
  regs__170 = _RAND_173[1:0];
  _RAND_174 = {1{`RANDOM}};
  regs__171 = _RAND_174[1:0];
  _RAND_175 = {1{`RANDOM}};
  regs__172 = _RAND_175[1:0];
  _RAND_176 = {1{`RANDOM}};
  regs__173 = _RAND_176[1:0];
  _RAND_177 = {1{`RANDOM}};
  regs__174 = _RAND_177[1:0];
  _RAND_178 = {1{`RANDOM}};
  regs__175 = _RAND_178[1:0];
  _RAND_179 = {1{`RANDOM}};
  regs__176 = _RAND_179[1:0];
  _RAND_180 = {1{`RANDOM}};
  regs__177 = _RAND_180[1:0];
  _RAND_181 = {1{`RANDOM}};
  regs__178 = _RAND_181[1:0];
  _RAND_182 = {1{`RANDOM}};
  regs__179 = _RAND_182[1:0];
  _RAND_183 = {1{`RANDOM}};
  regs__180 = _RAND_183[1:0];
  _RAND_184 = {1{`RANDOM}};
  regs__181 = _RAND_184[1:0];
  _RAND_185 = {1{`RANDOM}};
  regs__182 = _RAND_185[1:0];
  _RAND_186 = {1{`RANDOM}};
  regs__183 = _RAND_186[1:0];
  _RAND_187 = {1{`RANDOM}};
  regs__184 = _RAND_187[1:0];
  _RAND_188 = {1{`RANDOM}};
  regs__185 = _RAND_188[1:0];
  _RAND_189 = {1{`RANDOM}};
  regs__186 = _RAND_189[1:0];
  _RAND_190 = {1{`RANDOM}};
  regs__187 = _RAND_190[1:0];
  _RAND_191 = {1{`RANDOM}};
  regs__188 = _RAND_191[1:0];
  _RAND_192 = {1{`RANDOM}};
  regs__189 = _RAND_192[1:0];
  _RAND_193 = {1{`RANDOM}};
  regs__190 = _RAND_193[1:0];
  _RAND_194 = {1{`RANDOM}};
  regs__191 = _RAND_194[1:0];
  _RAND_195 = {1{`RANDOM}};
  regs__192 = _RAND_195[1:0];
  _RAND_196 = {1{`RANDOM}};
  regs__193 = _RAND_196[1:0];
  _RAND_197 = {1{`RANDOM}};
  regs__194 = _RAND_197[1:0];
  _RAND_198 = {1{`RANDOM}};
  regs__195 = _RAND_198[1:0];
  _RAND_199 = {1{`RANDOM}};
  regs__196 = _RAND_199[1:0];
  _RAND_200 = {1{`RANDOM}};
  regs__197 = _RAND_200[1:0];
  _RAND_201 = {1{`RANDOM}};
  regs__198 = _RAND_201[1:0];
  _RAND_202 = {1{`RANDOM}};
  regs__199 = _RAND_202[1:0];
  _RAND_203 = {1{`RANDOM}};
  regs__200 = _RAND_203[1:0];
  _RAND_204 = {1{`RANDOM}};
  regs__201 = _RAND_204[1:0];
  _RAND_205 = {1{`RANDOM}};
  regs__202 = _RAND_205[1:0];
  _RAND_206 = {1{`RANDOM}};
  regs__203 = _RAND_206[1:0];
  _RAND_207 = {1{`RANDOM}};
  regs__204 = _RAND_207[1:0];
  _RAND_208 = {1{`RANDOM}};
  regs__205 = _RAND_208[1:0];
  _RAND_209 = {1{`RANDOM}};
  regs__206 = _RAND_209[1:0];
  _RAND_210 = {1{`RANDOM}};
  regs__207 = _RAND_210[1:0];
  _RAND_211 = {1{`RANDOM}};
  regs__208 = _RAND_211[1:0];
  _RAND_212 = {1{`RANDOM}};
  regs__209 = _RAND_212[1:0];
  _RAND_213 = {1{`RANDOM}};
  regs__210 = _RAND_213[1:0];
  _RAND_214 = {1{`RANDOM}};
  regs__211 = _RAND_214[1:0];
  _RAND_215 = {1{`RANDOM}};
  regs__212 = _RAND_215[1:0];
  _RAND_216 = {1{`RANDOM}};
  regs__213 = _RAND_216[1:0];
  _RAND_217 = {1{`RANDOM}};
  regs__214 = _RAND_217[1:0];
  _RAND_218 = {1{`RANDOM}};
  regs__215 = _RAND_218[1:0];
  _RAND_219 = {1{`RANDOM}};
  regs__216 = _RAND_219[1:0];
  _RAND_220 = {1{`RANDOM}};
  regs__217 = _RAND_220[1:0];
  _RAND_221 = {1{`RANDOM}};
  regs__218 = _RAND_221[1:0];
  _RAND_222 = {1{`RANDOM}};
  regs__219 = _RAND_222[1:0];
  _RAND_223 = {1{`RANDOM}};
  regs__220 = _RAND_223[1:0];
  _RAND_224 = {1{`RANDOM}};
  regs__221 = _RAND_224[1:0];
  _RAND_225 = {1{`RANDOM}};
  regs__222 = _RAND_225[1:0];
  _RAND_226 = {1{`RANDOM}};
  regs__223 = _RAND_226[1:0];
  _RAND_227 = {1{`RANDOM}};
  regs__224 = _RAND_227[1:0];
  _RAND_228 = {1{`RANDOM}};
  regs__225 = _RAND_228[1:0];
  _RAND_229 = {1{`RANDOM}};
  regs__226 = _RAND_229[1:0];
  _RAND_230 = {1{`RANDOM}};
  regs__227 = _RAND_230[1:0];
  _RAND_231 = {1{`RANDOM}};
  regs__228 = _RAND_231[1:0];
  _RAND_232 = {1{`RANDOM}};
  regs__229 = _RAND_232[1:0];
  _RAND_233 = {1{`RANDOM}};
  regs__230 = _RAND_233[1:0];
  _RAND_234 = {1{`RANDOM}};
  regs__231 = _RAND_234[1:0];
  _RAND_235 = {1{`RANDOM}};
  regs__232 = _RAND_235[1:0];
  _RAND_236 = {1{`RANDOM}};
  regs__233 = _RAND_236[1:0];
  _RAND_237 = {1{`RANDOM}};
  regs__234 = _RAND_237[1:0];
  _RAND_238 = {1{`RANDOM}};
  regs__235 = _RAND_238[1:0];
  _RAND_239 = {1{`RANDOM}};
  regs__236 = _RAND_239[1:0];
  _RAND_240 = {1{`RANDOM}};
  regs__237 = _RAND_240[1:0];
  _RAND_241 = {1{`RANDOM}};
  regs__238 = _RAND_241[1:0];
  _RAND_242 = {1{`RANDOM}};
  regs__239 = _RAND_242[1:0];
  _RAND_243 = {1{`RANDOM}};
  regs__240 = _RAND_243[1:0];
  _RAND_244 = {1{`RANDOM}};
  regs__241 = _RAND_244[1:0];
  _RAND_245 = {1{`RANDOM}};
  regs__242 = _RAND_245[1:0];
  _RAND_246 = {1{`RANDOM}};
  regs__243 = _RAND_246[1:0];
  _RAND_247 = {1{`RANDOM}};
  regs__244 = _RAND_247[1:0];
  _RAND_248 = {1{`RANDOM}};
  regs__245 = _RAND_248[1:0];
  _RAND_249 = {1{`RANDOM}};
  regs__246 = _RAND_249[1:0];
  _RAND_250 = {1{`RANDOM}};
  regs__247 = _RAND_250[1:0];
  _RAND_251 = {1{`RANDOM}};
  regs__248 = _RAND_251[1:0];
  _RAND_252 = {1{`RANDOM}};
  regs__249 = _RAND_252[1:0];
  _RAND_253 = {1{`RANDOM}};
  regs__250 = _RAND_253[1:0];
  _RAND_254 = {1{`RANDOM}};
  regs__251 = _RAND_254[1:0];
  _RAND_255 = {1{`RANDOM}};
  regs__252 = _RAND_255[1:0];
  _RAND_256 = {1{`RANDOM}};
  regs__253 = _RAND_256[1:0];
  _RAND_257 = {1{`RANDOM}};
  regs__254 = _RAND_257[1:0];
  _RAND_258 = {1{`RANDOM}};
  regs__255 = _RAND_258[1:0];
  _RAND_259 = {1{`RANDOM}};
  regs__256 = _RAND_259[1:0];
  _RAND_260 = {1{`RANDOM}};
  regs__257 = _RAND_260[1:0];
  _RAND_261 = {1{`RANDOM}};
  regs__258 = _RAND_261[1:0];
  _RAND_262 = {1{`RANDOM}};
  regs__259 = _RAND_262[1:0];
  _RAND_263 = {1{`RANDOM}};
  regs__260 = _RAND_263[1:0];
  _RAND_264 = {1{`RANDOM}};
  regs__261 = _RAND_264[1:0];
  _RAND_265 = {1{`RANDOM}};
  regs__262 = _RAND_265[1:0];
  _RAND_266 = {1{`RANDOM}};
  regs__263 = _RAND_266[1:0];
  _RAND_267 = {1{`RANDOM}};
  regs__264 = _RAND_267[1:0];
  _RAND_268 = {1{`RANDOM}};
  regs__265 = _RAND_268[1:0];
  _RAND_269 = {1{`RANDOM}};
  regs__266 = _RAND_269[1:0];
  _RAND_270 = {1{`RANDOM}};
  regs__267 = _RAND_270[1:0];
  _RAND_271 = {1{`RANDOM}};
  regs__268 = _RAND_271[1:0];
  _RAND_272 = {1{`RANDOM}};
  regs__269 = _RAND_272[1:0];
  _RAND_273 = {1{`RANDOM}};
  regs__270 = _RAND_273[1:0];
  _RAND_274 = {1{`RANDOM}};
  regs__271 = _RAND_274[1:0];
  _RAND_275 = {1{`RANDOM}};
  regs__272 = _RAND_275[1:0];
  _RAND_276 = {1{`RANDOM}};
  regs__273 = _RAND_276[1:0];
  _RAND_277 = {1{`RANDOM}};
  regs__274 = _RAND_277[1:0];
  _RAND_278 = {1{`RANDOM}};
  regs__275 = _RAND_278[1:0];
  _RAND_279 = {1{`RANDOM}};
  regs__276 = _RAND_279[1:0];
  _RAND_280 = {1{`RANDOM}};
  regs__277 = _RAND_280[1:0];
  _RAND_281 = {1{`RANDOM}};
  regs__278 = _RAND_281[1:0];
  _RAND_282 = {1{`RANDOM}};
  regs__279 = _RAND_282[1:0];
  _RAND_283 = {1{`RANDOM}};
  regs__280 = _RAND_283[1:0];
  _RAND_284 = {1{`RANDOM}};
  regs__281 = _RAND_284[1:0];
  _RAND_285 = {1{`RANDOM}};
  regs__282 = _RAND_285[1:0];
  _RAND_286 = {1{`RANDOM}};
  regs__283 = _RAND_286[1:0];
  _RAND_287 = {1{`RANDOM}};
  regs__284 = _RAND_287[1:0];
  _RAND_288 = {1{`RANDOM}};
  regs__285 = _RAND_288[1:0];
  _RAND_289 = {1{`RANDOM}};
  regs__286 = _RAND_289[1:0];
  _RAND_290 = {1{`RANDOM}};
  regs__287 = _RAND_290[1:0];
  _RAND_291 = {1{`RANDOM}};
  regs__288 = _RAND_291[1:0];
  _RAND_292 = {1{`RANDOM}};
  regs__289 = _RAND_292[1:0];
  _RAND_293 = {1{`RANDOM}};
  regs__290 = _RAND_293[1:0];
  _RAND_294 = {1{`RANDOM}};
  regs__291 = _RAND_294[1:0];
  _RAND_295 = {1{`RANDOM}};
  regs__292 = _RAND_295[1:0];
  _RAND_296 = {1{`RANDOM}};
  regs__293 = _RAND_296[1:0];
  _RAND_297 = {1{`RANDOM}};
  regs__294 = _RAND_297[1:0];
  _RAND_298 = {1{`RANDOM}};
  regs__295 = _RAND_298[1:0];
  _RAND_299 = {1{`RANDOM}};
  regs__296 = _RAND_299[1:0];
  _RAND_300 = {1{`RANDOM}};
  regs__297 = _RAND_300[1:0];
  _RAND_301 = {1{`RANDOM}};
  regs__298 = _RAND_301[1:0];
  _RAND_302 = {1{`RANDOM}};
  regs__299 = _RAND_302[1:0];
  _RAND_303 = {1{`RANDOM}};
  regs__300 = _RAND_303[1:0];
  _RAND_304 = {1{`RANDOM}};
  regs__301 = _RAND_304[1:0];
  _RAND_305 = {1{`RANDOM}};
  regs__302 = _RAND_305[1:0];
  _RAND_306 = {1{`RANDOM}};
  regs__303 = _RAND_306[1:0];
  _RAND_307 = {1{`RANDOM}};
  regs__304 = _RAND_307[1:0];
  _RAND_308 = {1{`RANDOM}};
  regs__305 = _RAND_308[1:0];
  _RAND_309 = {1{`RANDOM}};
  regs__306 = _RAND_309[1:0];
  _RAND_310 = {1{`RANDOM}};
  regs__307 = _RAND_310[1:0];
  _RAND_311 = {1{`RANDOM}};
  regs__308 = _RAND_311[1:0];
  _RAND_312 = {1{`RANDOM}};
  regs__309 = _RAND_312[1:0];
  _RAND_313 = {1{`RANDOM}};
  regs__310 = _RAND_313[1:0];
  _RAND_314 = {1{`RANDOM}};
  regs__311 = _RAND_314[1:0];
  _RAND_315 = {1{`RANDOM}};
  regs__312 = _RAND_315[1:0];
  _RAND_316 = {1{`RANDOM}};
  regs__313 = _RAND_316[1:0];
  _RAND_317 = {1{`RANDOM}};
  regs__314 = _RAND_317[1:0];
  _RAND_318 = {1{`RANDOM}};
  regs__315 = _RAND_318[1:0];
  _RAND_319 = {1{`RANDOM}};
  regs__316 = _RAND_319[1:0];
  _RAND_320 = {1{`RANDOM}};
  regs__317 = _RAND_320[1:0];
  _RAND_321 = {1{`RANDOM}};
  regs__318 = _RAND_321[1:0];
  _RAND_322 = {1{`RANDOM}};
  regs__319 = _RAND_322[1:0];
  _RAND_323 = {1{`RANDOM}};
  regs__320 = _RAND_323[1:0];
  _RAND_324 = {1{`RANDOM}};
  regs__321 = _RAND_324[1:0];
  _RAND_325 = {1{`RANDOM}};
  regs__322 = _RAND_325[1:0];
  _RAND_326 = {1{`RANDOM}};
  regs__323 = _RAND_326[1:0];
  _RAND_327 = {1{`RANDOM}};
  regs__324 = _RAND_327[1:0];
  _RAND_328 = {1{`RANDOM}};
  regs__325 = _RAND_328[1:0];
  _RAND_329 = {1{`RANDOM}};
  regs__326 = _RAND_329[1:0];
  _RAND_330 = {1{`RANDOM}};
  regs__327 = _RAND_330[1:0];
  _RAND_331 = {1{`RANDOM}};
  regs__328 = _RAND_331[1:0];
  _RAND_332 = {1{`RANDOM}};
  regs__329 = _RAND_332[1:0];
  _RAND_333 = {1{`RANDOM}};
  regs__330 = _RAND_333[1:0];
  _RAND_334 = {1{`RANDOM}};
  regs__331 = _RAND_334[1:0];
  _RAND_335 = {1{`RANDOM}};
  regs__332 = _RAND_335[1:0];
  _RAND_336 = {1{`RANDOM}};
  regs__333 = _RAND_336[1:0];
  _RAND_337 = {1{`RANDOM}};
  regs__334 = _RAND_337[1:0];
  _RAND_338 = {1{`RANDOM}};
  regs__335 = _RAND_338[1:0];
  _RAND_339 = {1{`RANDOM}};
  regs__336 = _RAND_339[1:0];
  _RAND_340 = {1{`RANDOM}};
  regs__337 = _RAND_340[1:0];
  _RAND_341 = {1{`RANDOM}};
  regs__338 = _RAND_341[1:0];
  _RAND_342 = {1{`RANDOM}};
  regs__339 = _RAND_342[1:0];
  _RAND_343 = {1{`RANDOM}};
  regs__340 = _RAND_343[1:0];
  _RAND_344 = {1{`RANDOM}};
  regs__341 = _RAND_344[1:0];
  _RAND_345 = {1{`RANDOM}};
  regs__342 = _RAND_345[1:0];
  _RAND_346 = {1{`RANDOM}};
  regs__343 = _RAND_346[1:0];
  _RAND_347 = {1{`RANDOM}};
  regs__344 = _RAND_347[1:0];
  _RAND_348 = {1{`RANDOM}};
  regs__345 = _RAND_348[1:0];
  _RAND_349 = {1{`RANDOM}};
  regs__346 = _RAND_349[1:0];
  _RAND_350 = {1{`RANDOM}};
  regs__347 = _RAND_350[1:0];
  _RAND_351 = {1{`RANDOM}};
  regs__348 = _RAND_351[1:0];
  _RAND_352 = {1{`RANDOM}};
  regs__349 = _RAND_352[1:0];
  _RAND_353 = {1{`RANDOM}};
  regs__350 = _RAND_353[1:0];
  _RAND_354 = {1{`RANDOM}};
  regs__351 = _RAND_354[1:0];
  _RAND_355 = {1{`RANDOM}};
  regs__352 = _RAND_355[1:0];
  _RAND_356 = {1{`RANDOM}};
  regs__353 = _RAND_356[1:0];
  _RAND_357 = {1{`RANDOM}};
  regs__354 = _RAND_357[1:0];
  _RAND_358 = {1{`RANDOM}};
  regs__355 = _RAND_358[1:0];
  _RAND_359 = {1{`RANDOM}};
  regs__356 = _RAND_359[1:0];
  _RAND_360 = {1{`RANDOM}};
  regs__357 = _RAND_360[1:0];
  _RAND_361 = {1{`RANDOM}};
  regs__358 = _RAND_361[1:0];
  _RAND_362 = {1{`RANDOM}};
  regs__359 = _RAND_362[1:0];
  _RAND_363 = {1{`RANDOM}};
  regs__360 = _RAND_363[1:0];
  _RAND_364 = {1{`RANDOM}};
  regs__361 = _RAND_364[1:0];
  _RAND_365 = {1{`RANDOM}};
  regs__362 = _RAND_365[1:0];
  _RAND_366 = {1{`RANDOM}};
  regs__363 = _RAND_366[1:0];
  _RAND_367 = {1{`RANDOM}};
  regs__364 = _RAND_367[1:0];
  _RAND_368 = {1{`RANDOM}};
  regs__365 = _RAND_368[1:0];
  _RAND_369 = {1{`RANDOM}};
  regs__366 = _RAND_369[1:0];
  _RAND_370 = {1{`RANDOM}};
  regs__367 = _RAND_370[1:0];
  _RAND_371 = {1{`RANDOM}};
  regs__368 = _RAND_371[1:0];
  _RAND_372 = {1{`RANDOM}};
  regs__369 = _RAND_372[1:0];
  _RAND_373 = {1{`RANDOM}};
  regs__370 = _RAND_373[1:0];
  _RAND_374 = {1{`RANDOM}};
  regs__371 = _RAND_374[1:0];
  _RAND_375 = {1{`RANDOM}};
  regs__372 = _RAND_375[1:0];
  _RAND_376 = {1{`RANDOM}};
  regs__373 = _RAND_376[1:0];
  _RAND_377 = {1{`RANDOM}};
  regs__374 = _RAND_377[1:0];
  _RAND_378 = {1{`RANDOM}};
  regs__375 = _RAND_378[1:0];
  _RAND_379 = {1{`RANDOM}};
  regs__376 = _RAND_379[1:0];
  _RAND_380 = {1{`RANDOM}};
  regs__377 = _RAND_380[1:0];
  _RAND_381 = {1{`RANDOM}};
  regs__378 = _RAND_381[1:0];
  _RAND_382 = {1{`RANDOM}};
  regs__379 = _RAND_382[1:0];
  _RAND_383 = {1{`RANDOM}};
  regs__380 = _RAND_383[1:0];
  _RAND_384 = {1{`RANDOM}};
  regs__381 = _RAND_384[1:0];
  _RAND_385 = {1{`RANDOM}};
  regs__382 = _RAND_385[1:0];
  _RAND_386 = {1{`RANDOM}};
  regs__383 = _RAND_386[1:0];
  _RAND_387 = {1{`RANDOM}};
  regs__384 = _RAND_387[1:0];
  _RAND_388 = {1{`RANDOM}};
  regs__385 = _RAND_388[1:0];
  _RAND_389 = {1{`RANDOM}};
  regs__386 = _RAND_389[1:0];
  _RAND_390 = {1{`RANDOM}};
  regs__387 = _RAND_390[1:0];
  _RAND_391 = {1{`RANDOM}};
  regs__388 = _RAND_391[1:0];
  _RAND_392 = {1{`RANDOM}};
  regs__389 = _RAND_392[1:0];
  _RAND_393 = {1{`RANDOM}};
  regs__390 = _RAND_393[1:0];
  _RAND_394 = {1{`RANDOM}};
  regs__391 = _RAND_394[1:0];
  _RAND_395 = {1{`RANDOM}};
  regs__392 = _RAND_395[1:0];
  _RAND_396 = {1{`RANDOM}};
  regs__393 = _RAND_396[1:0];
  _RAND_397 = {1{`RANDOM}};
  regs__394 = _RAND_397[1:0];
  _RAND_398 = {1{`RANDOM}};
  regs__395 = _RAND_398[1:0];
  _RAND_399 = {1{`RANDOM}};
  regs__396 = _RAND_399[1:0];
  _RAND_400 = {1{`RANDOM}};
  regs__397 = _RAND_400[1:0];
  _RAND_401 = {1{`RANDOM}};
  regs__398 = _RAND_401[1:0];
  _RAND_402 = {1{`RANDOM}};
  regs__399 = _RAND_402[1:0];
  _RAND_403 = {1{`RANDOM}};
  regs__400 = _RAND_403[1:0];
  _RAND_404 = {1{`RANDOM}};
  regs__401 = _RAND_404[1:0];
  _RAND_405 = {1{`RANDOM}};
  regs__402 = _RAND_405[1:0];
  _RAND_406 = {1{`RANDOM}};
  regs__403 = _RAND_406[1:0];
  _RAND_407 = {1{`RANDOM}};
  regs__404 = _RAND_407[1:0];
  _RAND_408 = {1{`RANDOM}};
  regs__405 = _RAND_408[1:0];
  _RAND_409 = {1{`RANDOM}};
  regs__406 = _RAND_409[1:0];
  _RAND_410 = {1{`RANDOM}};
  regs__407 = _RAND_410[1:0];
  _RAND_411 = {1{`RANDOM}};
  regs__408 = _RAND_411[1:0];
  _RAND_412 = {1{`RANDOM}};
  regs__409 = _RAND_412[1:0];
  _RAND_413 = {1{`RANDOM}};
  regs__410 = _RAND_413[1:0];
  _RAND_414 = {1{`RANDOM}};
  regs__411 = _RAND_414[1:0];
  _RAND_415 = {1{`RANDOM}};
  regs__412 = _RAND_415[1:0];
  _RAND_416 = {1{`RANDOM}};
  regs__413 = _RAND_416[1:0];
  _RAND_417 = {1{`RANDOM}};
  regs__414 = _RAND_417[1:0];
  _RAND_418 = {1{`RANDOM}};
  regs__415 = _RAND_418[1:0];
  _RAND_419 = {1{`RANDOM}};
  regs__416 = _RAND_419[1:0];
  _RAND_420 = {1{`RANDOM}};
  regs__417 = _RAND_420[1:0];
  _RAND_421 = {1{`RANDOM}};
  regs__418 = _RAND_421[1:0];
  _RAND_422 = {1{`RANDOM}};
  regs__419 = _RAND_422[1:0];
  _RAND_423 = {1{`RANDOM}};
  regs__420 = _RAND_423[1:0];
  _RAND_424 = {1{`RANDOM}};
  regs__421 = _RAND_424[1:0];
  _RAND_425 = {1{`RANDOM}};
  regs__422 = _RAND_425[1:0];
  _RAND_426 = {1{`RANDOM}};
  regs__423 = _RAND_426[1:0];
  _RAND_427 = {1{`RANDOM}};
  regs__424 = _RAND_427[1:0];
  _RAND_428 = {1{`RANDOM}};
  regs__425 = _RAND_428[1:0];
  _RAND_429 = {1{`RANDOM}};
  regs__426 = _RAND_429[1:0];
  _RAND_430 = {1{`RANDOM}};
  regs__427 = _RAND_430[1:0];
  _RAND_431 = {1{`RANDOM}};
  regs__428 = _RAND_431[1:0];
  _RAND_432 = {1{`RANDOM}};
  regs__429 = _RAND_432[1:0];
  _RAND_433 = {1{`RANDOM}};
  regs__430 = _RAND_433[1:0];
  _RAND_434 = {1{`RANDOM}};
  regs__431 = _RAND_434[1:0];
  _RAND_435 = {1{`RANDOM}};
  regs__432 = _RAND_435[1:0];
  _RAND_436 = {1{`RANDOM}};
  regs__433 = _RAND_436[1:0];
  _RAND_437 = {1{`RANDOM}};
  regs__434 = _RAND_437[1:0];
  _RAND_438 = {1{`RANDOM}};
  regs__435 = _RAND_438[1:0];
  _RAND_439 = {1{`RANDOM}};
  regs__436 = _RAND_439[1:0];
  _RAND_440 = {1{`RANDOM}};
  regs__437 = _RAND_440[1:0];
  _RAND_441 = {1{`RANDOM}};
  regs__438 = _RAND_441[1:0];
  _RAND_442 = {1{`RANDOM}};
  regs__439 = _RAND_442[1:0];
  _RAND_443 = {1{`RANDOM}};
  regs__440 = _RAND_443[1:0];
  _RAND_444 = {1{`RANDOM}};
  regs__441 = _RAND_444[1:0];
  _RAND_445 = {1{`RANDOM}};
  regs__442 = _RAND_445[1:0];
  _RAND_446 = {1{`RANDOM}};
  regs__443 = _RAND_446[1:0];
  _RAND_447 = {1{`RANDOM}};
  regs__444 = _RAND_447[1:0];
  _RAND_448 = {1{`RANDOM}};
  regs__445 = _RAND_448[1:0];
  _RAND_449 = {1{`RANDOM}};
  regs__446 = _RAND_449[1:0];
  _RAND_450 = {1{`RANDOM}};
  regs__447 = _RAND_450[1:0];
  _RAND_451 = {1{`RANDOM}};
  regs__448 = _RAND_451[1:0];
  _RAND_452 = {1{`RANDOM}};
  regs__449 = _RAND_452[1:0];
  _RAND_453 = {1{`RANDOM}};
  regs__450 = _RAND_453[1:0];
  _RAND_454 = {1{`RANDOM}};
  regs__451 = _RAND_454[1:0];
  _RAND_455 = {1{`RANDOM}};
  regs__452 = _RAND_455[1:0];
  _RAND_456 = {1{`RANDOM}};
  regs__453 = _RAND_456[1:0];
  _RAND_457 = {1{`RANDOM}};
  regs__454 = _RAND_457[1:0];
  _RAND_458 = {1{`RANDOM}};
  regs__455 = _RAND_458[1:0];
  _RAND_459 = {1{`RANDOM}};
  regs__456 = _RAND_459[1:0];
  _RAND_460 = {1{`RANDOM}};
  regs__457 = _RAND_460[1:0];
  _RAND_461 = {1{`RANDOM}};
  regs__458 = _RAND_461[1:0];
  _RAND_462 = {1{`RANDOM}};
  regs__459 = _RAND_462[1:0];
  _RAND_463 = {1{`RANDOM}};
  regs__460 = _RAND_463[1:0];
  _RAND_464 = {1{`RANDOM}};
  regs__461 = _RAND_464[1:0];
  _RAND_465 = {1{`RANDOM}};
  regs__462 = _RAND_465[1:0];
  _RAND_466 = {1{`RANDOM}};
  regs__463 = _RAND_466[1:0];
  _RAND_467 = {1{`RANDOM}};
  regs__464 = _RAND_467[1:0];
  _RAND_468 = {1{`RANDOM}};
  regs__465 = _RAND_468[1:0];
  _RAND_469 = {1{`RANDOM}};
  regs__466 = _RAND_469[1:0];
  _RAND_470 = {1{`RANDOM}};
  regs__467 = _RAND_470[1:0];
  _RAND_471 = {1{`RANDOM}};
  regs__468 = _RAND_471[1:0];
  _RAND_472 = {1{`RANDOM}};
  regs__469 = _RAND_472[1:0];
  _RAND_473 = {1{`RANDOM}};
  regs__470 = _RAND_473[1:0];
  _RAND_474 = {1{`RANDOM}};
  regs__471 = _RAND_474[1:0];
  _RAND_475 = {1{`RANDOM}};
  regs__472 = _RAND_475[1:0];
  _RAND_476 = {1{`RANDOM}};
  regs__473 = _RAND_476[1:0];
  _RAND_477 = {1{`RANDOM}};
  regs__474 = _RAND_477[1:0];
  _RAND_478 = {1{`RANDOM}};
  regs__475 = _RAND_478[1:0];
  _RAND_479 = {1{`RANDOM}};
  regs__476 = _RAND_479[1:0];
  _RAND_480 = {1{`RANDOM}};
  regs__477 = _RAND_480[1:0];
  _RAND_481 = {1{`RANDOM}};
  regs__478 = _RAND_481[1:0];
  _RAND_482 = {1{`RANDOM}};
  regs__479 = _RAND_482[1:0];
  _RAND_483 = {1{`RANDOM}};
  regs__480 = _RAND_483[1:0];
  _RAND_484 = {1{`RANDOM}};
  regs__481 = _RAND_484[1:0];
  _RAND_485 = {1{`RANDOM}};
  regs__482 = _RAND_485[1:0];
  _RAND_486 = {1{`RANDOM}};
  regs__483 = _RAND_486[1:0];
  _RAND_487 = {1{`RANDOM}};
  regs__484 = _RAND_487[1:0];
  _RAND_488 = {1{`RANDOM}};
  regs__485 = _RAND_488[1:0];
  _RAND_489 = {1{`RANDOM}};
  regs__486 = _RAND_489[1:0];
  _RAND_490 = {1{`RANDOM}};
  regs__487 = _RAND_490[1:0];
  _RAND_491 = {1{`RANDOM}};
  regs__488 = _RAND_491[1:0];
  _RAND_492 = {1{`RANDOM}};
  regs__489 = _RAND_492[1:0];
  _RAND_493 = {1{`RANDOM}};
  regs__490 = _RAND_493[1:0];
  _RAND_494 = {1{`RANDOM}};
  regs__491 = _RAND_494[1:0];
  _RAND_495 = {1{`RANDOM}};
  regs__492 = _RAND_495[1:0];
  _RAND_496 = {1{`RANDOM}};
  regs__493 = _RAND_496[1:0];
  _RAND_497 = {1{`RANDOM}};
  regs__494 = _RAND_497[1:0];
  _RAND_498 = {1{`RANDOM}};
  regs__495 = _RAND_498[1:0];
  _RAND_499 = {1{`RANDOM}};
  regs__496 = _RAND_499[1:0];
  _RAND_500 = {1{`RANDOM}};
  regs__497 = _RAND_500[1:0];
  _RAND_501 = {1{`RANDOM}};
  regs__498 = _RAND_501[1:0];
  _RAND_502 = {1{`RANDOM}};
  regs__499 = _RAND_502[1:0];
  _RAND_503 = {1{`RANDOM}};
  regs__500 = _RAND_503[1:0];
  _RAND_504 = {1{`RANDOM}};
  regs__501 = _RAND_504[1:0];
  _RAND_505 = {1{`RANDOM}};
  regs__502 = _RAND_505[1:0];
  _RAND_506 = {1{`RANDOM}};
  regs__503 = _RAND_506[1:0];
  _RAND_507 = {1{`RANDOM}};
  regs__504 = _RAND_507[1:0];
  _RAND_508 = {1{`RANDOM}};
  regs__505 = _RAND_508[1:0];
  _RAND_509 = {1{`RANDOM}};
  regs__506 = _RAND_509[1:0];
  _RAND_510 = {1{`RANDOM}};
  regs__507 = _RAND_510[1:0];
  _RAND_511 = {1{`RANDOM}};
  regs__508 = _RAND_511[1:0];
  _RAND_512 = {1{`RANDOM}};
  regs__509 = _RAND_512[1:0];
  _RAND_513 = {1{`RANDOM}};
  regs__510 = _RAND_513[1:0];
  _RAND_514 = {1{`RANDOM}};
  regs__511 = _RAND_514[1:0];
  _RAND_515 = {1{`RANDOM}};
  phtTaken = _RAND_515[0:0];
  _RAND_516 = {2{`RANDOM}};
  regs_1_0 = _RAND_516[38:0];
  _RAND_517 = {2{`RANDOM}};
  regs_1_1 = _RAND_517[38:0];
  _RAND_518 = {2{`RANDOM}};
  regs_1_2 = _RAND_518[38:0];
  _RAND_519 = {2{`RANDOM}};
  regs_1_3 = _RAND_519[38:0];
  _RAND_520 = {2{`RANDOM}};
  regs_1_4 = _RAND_520[38:0];
  _RAND_521 = {2{`RANDOM}};
  regs_1_5 = _RAND_521[38:0];
  _RAND_522 = {2{`RANDOM}};
  regs_1_6 = _RAND_522[38:0];
  _RAND_523 = {2{`RANDOM}};
  regs_1_7 = _RAND_523[38:0];
  _RAND_524 = {2{`RANDOM}};
  regs_1_8 = _RAND_524[38:0];
  _RAND_525 = {2{`RANDOM}};
  regs_1_9 = _RAND_525[38:0];
  _RAND_526 = {2{`RANDOM}};
  regs_1_10 = _RAND_526[38:0];
  _RAND_527 = {2{`RANDOM}};
  regs_1_11 = _RAND_527[38:0];
  _RAND_528 = {2{`RANDOM}};
  regs_1_12 = _RAND_528[38:0];
  _RAND_529 = {2{`RANDOM}};
  regs_1_13 = _RAND_529[38:0];
  _RAND_530 = {2{`RANDOM}};
  regs_1_14 = _RAND_530[38:0];
  _RAND_531 = {2{`RANDOM}};
  regs_1_15 = _RAND_531[38:0];
  _RAND_532 = {1{`RANDOM}};
  sp_value = _RAND_532[3:0];
  _RAND_533 = {2{`RANDOM}};
  rasTarget = _RAND_533[38:0];
  _RAND_534 = {1{`RANDOM}};
  cnt = _RAND_534[1:0];
  _RAND_535 = {1{`RANDOM}};
  reqLatch_valid = _RAND_535[0:0];
  _RAND_536 = {2{`RANDOM}};
  reqLatch_pc = _RAND_536[38:0];
  _RAND_537 = {1{`RANDOM}};
  reqLatch_actualTaken = _RAND_537[0:0];
  _RAND_538 = {1{`RANDOM}};
  reqLatch_fuOpType = _RAND_538[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IFU_inorder(
  input         clock,
  input         reset,
  input         io_imem_req_ready, // @[src/main/scala/nutcore/frontend/IFU.scala 329:14]
  output        io_imem_req_valid, // @[src/main/scala/nutcore/frontend/IFU.scala 329:14]
  output [38:0] io_imem_req_bits_addr, // @[src/main/scala/nutcore/frontend/IFU.scala 329:14]
  output [81:0] io_imem_req_bits_user, // @[src/main/scala/nutcore/frontend/IFU.scala 329:14]
  output        io_imem_resp_ready, // @[src/main/scala/nutcore/frontend/IFU.scala 329:14]
  input         io_imem_resp_valid, // @[src/main/scala/nutcore/frontend/IFU.scala 329:14]
  input  [63:0] io_imem_resp_bits_rdata, // @[src/main/scala/nutcore/frontend/IFU.scala 329:14]
  input  [81:0] io_imem_resp_bits_user, // @[src/main/scala/nutcore/frontend/IFU.scala 329:14]
  input         io_out_ready, // @[src/main/scala/nutcore/frontend/IFU.scala 329:14]
  output        io_out_valid, // @[src/main/scala/nutcore/frontend/IFU.scala 329:14]
  output [63:0] io_out_bits_instr, // @[src/main/scala/nutcore/frontend/IFU.scala 329:14]
  output [38:0] io_out_bits_pc, // @[src/main/scala/nutcore/frontend/IFU.scala 329:14]
  output [38:0] io_out_bits_pnpc, // @[src/main/scala/nutcore/frontend/IFU.scala 329:14]
  output [3:0]  io_out_bits_brIdx, // @[src/main/scala/nutcore/frontend/IFU.scala 329:14]
  input  [38:0] io_redirect_target, // @[src/main/scala/nutcore/frontend/IFU.scala 329:14]
  input         io_redirect_valid, // @[src/main/scala/nutcore/frontend/IFU.scala 329:14]
  output [3:0]  io_flushVec, // @[src/main/scala/nutcore/frontend/IFU.scala 329:14]
  input         flushICache,
  input         REG_valid,
  input  [38:0] REG_pc,
  input         REG_isMissPredict,
  input  [38:0] REG_actualTarget,
  input         REG_actualTaken,
  input  [6:0]  REG_fuOpType,
  input  [1:0]  REG_btbType,
  input         REG_isRVC,
  input         flushTLB
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  bp1_clock; // @[src/main/scala/nutcore/frontend/IFU.scala 345:19]
  wire  bp1_reset; // @[src/main/scala/nutcore/frontend/IFU.scala 345:19]
  wire  bp1_io_in_pc_valid; // @[src/main/scala/nutcore/frontend/IFU.scala 345:19]
  wire [38:0] bp1_io_in_pc_bits; // @[src/main/scala/nutcore/frontend/IFU.scala 345:19]
  wire [38:0] bp1_io_out_target; // @[src/main/scala/nutcore/frontend/IFU.scala 345:19]
  wire  bp1_io_out_valid; // @[src/main/scala/nutcore/frontend/IFU.scala 345:19]
  wire  bp1_io_flush; // @[src/main/scala/nutcore/frontend/IFU.scala 345:19]
  wire [2:0] bp1_io_brIdx; // @[src/main/scala/nutcore/frontend/IFU.scala 345:19]
  wire  bp1_io_crosslineJump; // @[src/main/scala/nutcore/frontend/IFU.scala 345:19]
  wire  bp1_MOUFlushICache; // @[src/main/scala/nutcore/frontend/IFU.scala 345:19]
  wire  bp1_bpuUpdateReq_valid; // @[src/main/scala/nutcore/frontend/IFU.scala 345:19]
  wire [38:0] bp1_bpuUpdateReq_pc; // @[src/main/scala/nutcore/frontend/IFU.scala 345:19]
  wire  bp1_bpuUpdateReq_isMissPredict; // @[src/main/scala/nutcore/frontend/IFU.scala 345:19]
  wire [38:0] bp1_bpuUpdateReq_actualTarget; // @[src/main/scala/nutcore/frontend/IFU.scala 345:19]
  wire  bp1_bpuUpdateReq_actualTaken; // @[src/main/scala/nutcore/frontend/IFU.scala 345:19]
  wire [6:0] bp1_bpuUpdateReq_fuOpType; // @[src/main/scala/nutcore/frontend/IFU.scala 345:19]
  wire [1:0] bp1_bpuUpdateReq_btbType; // @[src/main/scala/nutcore/frontend/IFU.scala 345:19]
  wire  bp1_bpuUpdateReq_isRVC; // @[src/main/scala/nutcore/frontend/IFU.scala 345:19]
  wire  bp1_MOUFlushTLB; // @[src/main/scala/nutcore/frontend/IFU.scala 345:19]
  reg [38:0] pc; // @[src/main/scala/nutcore/frontend/IFU.scala 341:19]
  wire  _pcUpdate_T = io_imem_req_ready & io_imem_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  pcUpdate = io_redirect_valid | _pcUpdate_T; // @[src/main/scala/nutcore/frontend/IFU.scala 342:36]
  wire [38:0] _snpc_T_2 = pc + 39'h2; // @[src/main/scala/nutcore/frontend/IFU.scala 343:28]
  wire [38:0] _snpc_T_4 = pc + 39'h4; // @[src/main/scala/nutcore/frontend/IFU.scala 343:38]
  wire [38:0] snpc = pc[1] ? _snpc_T_2 : _snpc_T_4; // @[src/main/scala/nutcore/frontend/IFU.scala 343:17]
  reg  crosslineJumpLatch; // @[src/main/scala/nutcore/frontend/IFU.scala 348:35]
  reg [38:0] crosslineJumpTarget; // @[src/main/scala/nutcore/frontend/IFU.scala 352:38]
  wire [38:0] pnpc = bp1_io_crosslineJump ? snpc : bp1_io_out_target; // @[src/main/scala/nutcore/frontend/IFU.scala 357:17]
  wire [38:0] _npc_T = bp1_io_out_valid ? pnpc : snpc; // @[src/main/scala/nutcore/frontend/IFU.scala 359:104]
  wire [38:0] _npc_T_1 = crosslineJumpLatch ? crosslineJumpTarget : _npc_T; // @[src/main/scala/nutcore/frontend/IFU.scala 359:59]
  wire [38:0] npc = io_redirect_valid ? io_redirect_target : _npc_T_1; // @[src/main/scala/nutcore/frontend/IFU.scala 359:16]
  wire  _npcIsSeq_T = bp1_io_out_valid ? 1'h0 : 1'h1; // @[src/main/scala/nutcore/frontend/IFU.scala 360:114]
  wire  _npcIsSeq_T_2 = crosslineJumpLatch ? 1'h0 : bp1_io_crosslineJump | _npcIsSeq_T; // @[src/main/scala/nutcore/frontend/IFU.scala 360:54]
  wire  npcIsSeq = io_redirect_valid ? 1'h0 : _npcIsSeq_T_2; // @[src/main/scala/nutcore/frontend/IFU.scala 360:21]
  wire [2:0] _brIdx_T = io_redirect_valid ? 3'h0 : bp1_io_brIdx; // @[src/main/scala/nutcore/frontend/IFU.scala 368:29]
  wire [42:0] x6_hi = {npcIsSeq,_brIdx_T,npc}; // @[src/main/scala/nutcore/frontend/IFU.scala 390:82]
  wire  _T_18 = io_imem_resp_ready & io_imem_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_3 = io_imem_req_valid | r; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  _T_19 = |io_flushVec; // @[src/main/scala/nutcore/frontend/IFU.scala 413:37]
  BPU_inorder bp1 ( // @[src/main/scala/nutcore/frontend/IFU.scala 345:19]
    .clock(bp1_clock),
    .reset(bp1_reset),
    .io_in_pc_valid(bp1_io_in_pc_valid),
    .io_in_pc_bits(bp1_io_in_pc_bits),
    .io_out_target(bp1_io_out_target),
    .io_out_valid(bp1_io_out_valid),
    .io_flush(bp1_io_flush),
    .io_brIdx(bp1_io_brIdx),
    .io_crosslineJump(bp1_io_crosslineJump),
    .MOUFlushICache(bp1_MOUFlushICache),
    .bpuUpdateReq_valid(bp1_bpuUpdateReq_valid),
    .bpuUpdateReq_pc(bp1_bpuUpdateReq_pc),
    .bpuUpdateReq_isMissPredict(bp1_bpuUpdateReq_isMissPredict),
    .bpuUpdateReq_actualTarget(bp1_bpuUpdateReq_actualTarget),
    .bpuUpdateReq_actualTaken(bp1_bpuUpdateReq_actualTaken),
    .bpuUpdateReq_fuOpType(bp1_bpuUpdateReq_fuOpType),
    .bpuUpdateReq_btbType(bp1_bpuUpdateReq_btbType),
    .bpuUpdateReq_isRVC(bp1_bpuUpdateReq_isRVC),
    .MOUFlushTLB(bp1_MOUFlushTLB)
  );
  assign io_imem_req_valid = io_out_ready; // @[src/main/scala/nutcore/frontend/IFU.scala 391:21]
  assign io_imem_req_bits_addr = {pc[38:1],1'h0}; // @[src/main/scala/nutcore/frontend/IFU.scala 389:36]
  assign io_imem_req_bits_user = {x6_hi,pc}; // @[src/main/scala/nutcore/frontend/IFU.scala 390:82]
  assign io_imem_resp_ready = io_out_ready | io_flushVec[0]; // @[src/main/scala/nutcore/frontend/IFU.scala 393:38]
  assign io_out_valid = io_imem_resp_valid & ~io_flushVec[0]; // @[src/main/scala/nutcore/frontend/IFU.scala 410:38]
  assign io_out_bits_instr = io_imem_resp_bits_rdata; // @[src/main/scala/nutcore/frontend/IFU.scala 403:21]
  assign io_out_bits_pc = io_imem_resp_bits_user[38:0]; // @[src/main/scala/nutcore/frontend/IFU.scala 405:24]
  assign io_out_bits_pnpc = io_imem_resp_bits_user[77:39]; // @[src/main/scala/nutcore/frontend/IFU.scala 406:26]
  assign io_out_bits_brIdx = io_imem_resp_bits_user[81:78]; // @[src/main/scala/nutcore/frontend/IFU.scala 407:27]
  assign io_flushVec = io_redirect_valid ? 4'hf : 4'h0; // @[src/main/scala/nutcore/frontend/IFU.scala 386:21]
  assign bp1_clock = clock;
  assign bp1_reset = reset;
  assign bp1_io_in_pc_valid = io_imem_req_ready & io_imem_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  assign bp1_io_in_pc_bits = io_redirect_valid ? io_redirect_target : _npc_T_1; // @[src/main/scala/nutcore/frontend/IFU.scala 359:16]
  assign bp1_io_flush = io_redirect_valid; // @[src/main/scala/nutcore/frontend/IFU.scala 377:16]
  assign bp1_MOUFlushICache = flushICache;
  assign bp1_bpuUpdateReq_valid = REG_valid;
  assign bp1_bpuUpdateReq_pc = REG_pc;
  assign bp1_bpuUpdateReq_isMissPredict = REG_isMissPredict;
  assign bp1_bpuUpdateReq_actualTarget = REG_actualTarget;
  assign bp1_bpuUpdateReq_actualTaken = REG_actualTaken;
  assign bp1_bpuUpdateReq_fuOpType = REG_fuOpType;
  assign bp1_bpuUpdateReq_btbType = REG_btbType;
  assign bp1_bpuUpdateReq_isRVC = REG_isRVC;
  assign bp1_MOUFlushTLB = flushTLB;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/frontend/IFU.scala 341:19]
      pc <= 39'h80000000; // @[src/main/scala/nutcore/frontend/IFU.scala 341:19]
    end else if (pcUpdate) begin // @[src/main/scala/nutcore/frontend/IFU.scala 379:19]
      if (io_redirect_valid) begin // @[src/main/scala/nutcore/frontend/IFU.scala 359:16]
        pc <= io_redirect_target;
      end else if (crosslineJumpLatch) begin // @[src/main/scala/nutcore/frontend/IFU.scala 359:59]
        pc <= crosslineJumpTarget;
      end else begin
        pc <= _npc_T;
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/frontend/IFU.scala 348:35]
      crosslineJumpLatch <= 1'h0; // @[src/main/scala/nutcore/frontend/IFU.scala 348:35]
    end else if (pcUpdate | bp1_io_flush) begin // @[src/main/scala/nutcore/frontend/IFU.scala 349:34]
      if (bp1_io_flush) begin // @[src/main/scala/nutcore/frontend/IFU.scala 350:30]
        crosslineJumpLatch <= 1'h0;
      end else begin
        crosslineJumpLatch <= bp1_io_crosslineJump & ~crosslineJumpLatch;
      end
    end
    if (bp1_io_crosslineJump) begin // @[src/main/scala/nutcore/frontend/IFU.scala 352:38]
      crosslineJumpTarget <= bp1_io_out_target; // @[src/main/scala/nutcore/frontend/IFU.scala 352:38]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (_T_18) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      r <= _GEN_3;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  pc = _RAND_0[38:0];
  _RAND_1 = {1{`RANDOM}};
  crosslineJumpLatch = _RAND_1[0:0];
  _RAND_2 = {2{`RANDOM}};
  crosslineJumpTarget = _RAND_2[38:0];
  _RAND_3 = {1{`RANDOM}};
  r = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module NaiveRVCAlignBuffer(
  input         clock,
  input         reset,
  output        io_in_ready, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_valid, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input  [63:0] io_in_bits_instr, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input  [38:0] io_in_bits_pc, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input  [38:0] io_in_bits_pnpc, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input  [3:0]  io_in_bits_brIdx, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_out_ready, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  output        io_out_valid, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  output [63:0] io_out_bits_instr, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  output [38:0] io_out_bits_pc, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  output [38:0] io_out_bits_pnpc, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  output [3:0]  io_out_bits_brIdx, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_flush // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 39:22]
  wire [79:0] instIn = {16'h0,io_in_bits_instr}; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 42:19]
  reg [15:0] specialInstR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:25]
  wire [31:0] _instr_T_4 = {instIn[15:0],specialInstR}; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 90:73]
  wire  _pcOffset_T = state == 2'h0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 41:28]
  reg [2:0] pcOffsetR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 40:26]
  wire [2:0] pcOffset = state == 2'h0 ? io_in_bits_pc[2:0] : pcOffsetR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 41:21]
  wire  _instr_T_9 = 3'h0 == pcOffset; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [31:0] _instr_T_13 = _instr_T_9 ? instIn[31:0] : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _instr_T_10 = 3'h2 == pcOffset; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [31:0] _instr_T_14 = _instr_T_10 ? instIn[47:16] : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _instr_T_17 = _instr_T_13 | _instr_T_14; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _instr_T_11 = 3'h4 == pcOffset; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [31:0] _instr_T_15 = _instr_T_11 ? instIn[63:32] : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _instr_T_18 = _instr_T_17 | _instr_T_15; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _instr_T_12 = 3'h6 == pcOffset; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [31:0] _instr_T_16 = _instr_T_12 ? instIn[79:48] : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _instr_T_19 = _instr_T_18 | _instr_T_16; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] instr = state == 2'h2 | state == 2'h3 ? _instr_T_4 : _instr_T_19; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 90:15]
  wire  isRVC = instr[1:0] != 2'h3; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 34:26]
  wire  _rvcFinish_T = pcOffset == 3'h0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 48:28]
  wire  _rvcFinish_T_1 = ~isRVC; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 48:40]
  wire  _rvcFinish_T_5 = pcOffset == 3'h4; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 48:72]
  wire  _rvcFinish_T_11 = pcOffset == 3'h2; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 48:116]
  wire  _rvcFinish_T_16 = pcOffset == 3'h6; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 48:159]
  wire  rvcFinish = pcOffset == 3'h0 & (~isRVC | io_in_bits_brIdx[0]) | pcOffset == 3'h4 & (~isRVC | io_in_bits_brIdx[0]
    ) | pcOffset == 3'h2 & (isRVC | io_in_bits_brIdx[1]) | pcOffset == 3'h6 & isRVC; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 48:147]
  wire  _rvcNext_T_13 = _rvcFinish_T_11 & _rvcFinish_T_1; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 51:122]
  wire  _rvcNext_T_15 = ~io_in_bits_brIdx[1]; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 51:135]
  wire  rvcNext = _rvcFinish_T & (isRVC & ~io_in_bits_brIdx[0]) | _rvcFinish_T_5 & (isRVC & ~io_in_bits_brIdx[0]) |
    _rvcFinish_T_11 & _rvcFinish_T_1 & ~io_in_bits_brIdx[1]; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 51:102]
  wire  _rvcSpecial_T_2 = _rvcFinish_T_16 & _rvcFinish_T_1; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 52:37]
  wire  rvcSpecial = _rvcFinish_T_16 & _rvcFinish_T_1 & ~io_in_bits_brIdx[2]; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 52:47]
  wire  rvcSpecialJump = _rvcSpecial_T_2 & io_in_bits_brIdx[2]; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 53:51]
  wire  pnpcIsSeq = io_in_bits_brIdx[3]; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 54:24]
  wire  _flushIFU_T_2 = _pcOffset_T | state == 2'h1; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 57:36]
  wire  flushIFU = (_pcOffset_T | state == 2'h1) & rvcSpecial & io_in_valid & ~pnpcIsSeq; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 57:87]
  wire  _T_2 = ~reset; // @[src/main/scala/utils/Debug.scala 56:24]
  wire  loadNextInstline = _flushIFU_T_2 & (rvcSpecial | rvcSpecialJump) & io_in_valid & pnpcIsSeq; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 60:115]
  reg [38:0] specialPCR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 64:23]
  reg [38:0] specialNPCR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 65:24]
  wire  rvcForceLoadNext = _rvcNext_T_13 & io_in_bits_pnpc[2:0] == 3'h4 & _rvcNext_T_15; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 69:86]
  wire  _canGo_T = rvcFinish | rvcNext; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 100:28]
  wire  _canIn_T = rvcFinish | rvcForceLoadNext; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:28]
  wire [38:0] _pnpcOut_T_1 = io_in_bits_pc + 39'h2; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 103:76]
  wire [38:0] _pnpcOut_T_3 = io_in_bits_pc + 39'h4; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 103:95]
  wire [38:0] _pnpcOut_T_4 = isRVC ? _pnpcOut_T_1 : _pnpcOut_T_3; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 103:55]
  wire [38:0] _pnpcOut_T_5 = rvcFinish ? io_in_bits_pnpc : _pnpcOut_T_4; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 103:23]
  wire  _T_11 = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [1:0] _GEN_0 = _T_11 & rvcFinish ? 2'h0 : state; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 104:{39,46} 39:22]
  wire [2:0] _pcOffsetR_T = isRVC ? 3'h2 : 3'h4; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 107:38]
  wire [2:0] _pcOffsetR_T_2 = pcOffset + _pcOffsetR_T; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 107:33]
  wire [1:0] _GEN_1 = _T_11 & rvcNext ? 2'h1 : _GEN_0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 105:37 106:17]
  wire [2:0] _GEN_2 = _T_11 & rvcNext ? _pcOffsetR_T_2 : pcOffsetR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 105:37 107:21 40:26]
  wire [1:0] _GEN_3 = rvcSpecial & io_in_valid ? 2'h2 : _GEN_1; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 109:40 110:17]
  wire [38:0] _pcOut_T_2 = {io_in_bits_pc[38:3],pcOffsetR}; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 126:21]
  wire [38:0] _GEN_27 = 2'h3 == state ? specialPCR : 39'h0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 161:15 98:18 62:23]
  wire [38:0] _GEN_32 = 2'h2 == state ? specialPCR : _GEN_27; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 149:15 98:18]
  wire [38:0] _GEN_40 = 2'h1 == state ? _pcOut_T_2 : _GEN_32; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 126:15 98:18]
  wire [38:0] pcOut = 2'h0 == state ? io_in_bits_pc : _GEN_40; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 102:15 98:18]
  wire [38:0] _GEN_4 = rvcSpecial & io_in_valid ? pcOut : specialPCR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 109:40 111:22 64:23]
  wire [15:0] _GEN_5 = rvcSpecial & io_in_valid ? io_in_bits_instr[63:48] : specialInstR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 109:40 112:24 66:25]
  wire [1:0] _GEN_7 = rvcSpecialJump & io_in_valid ? 2'h3 : _GEN_3; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 115:44 116:17]
  wire [38:0] _GEN_8 = rvcSpecialJump & io_in_valid ? pcOut : _GEN_4; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 115:44 117:22]
  wire [38:0] _GEN_9 = rvcSpecialJump & io_in_valid ? io_in_bits_pnpc : specialNPCR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 115:44 118:23 65:24]
  wire [15:0] _GEN_10 = rvcSpecialJump & io_in_valid ? io_in_bits_instr[63:48] : _GEN_5; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 115:44 119:24]
  wire [38:0] _pnpcOut_T_7 = pcOut + 39'h2; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 127:68]
  wire [38:0] _pnpcOut_T_9 = pcOut + 39'h4; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 127:79]
  wire [38:0] _pnpcOut_T_10 = isRVC ? _pnpcOut_T_7 : _pnpcOut_T_9; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 127:55]
  wire [38:0] _pnpcOut_T_11 = rvcFinish ? io_in_bits_pnpc : _pnpcOut_T_10; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 127:23]
  wire [38:0] _pnpcOut_T_13 = specialPCR + 39'h4; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 150:31]
  wire [1:0] _GEN_24 = _T_11 ? 2'h1 : state; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 154:26 155:17 39:22]
  wire [2:0] _GEN_25 = _T_11 ? 3'h2 : pcOffsetR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 154:26 156:21 40:26]
  wire [1:0] _GEN_26 = _T_11 ? 2'h0 : state; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 166:26 167:17 39:22]
  wire [38:0] _GEN_28 = 2'h3 == state ? specialNPCR : 39'h0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 162:17 98:18 63:25]
  wire  _GEN_29 = 2'h3 == state & io_in_valid; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 164:15 98:18 44:23]
  wire [1:0] _GEN_31 = 2'h3 == state ? _GEN_26 : state; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 98:18 39:22]
  wire [38:0] _GEN_33 = 2'h2 == state ? _pnpcOut_T_13 : _GEN_28; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 150:17 98:18]
  wire  _GEN_34 = 2'h2 == state ? io_in_valid : _GEN_29; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 152:15 98:18]
  wire  _GEN_35 = 2'h2 == state ? 1'h0 : 2'h3 == state; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 153:15 98:18]
  wire [1:0] _GEN_36 = 2'h2 == state ? _GEN_24 : _GEN_31; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 98:18]
  wire [2:0] _GEN_37 = 2'h2 == state ? _GEN_25 : pcOffsetR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 98:18 40:26]
  wire  _GEN_38 = 2'h1 == state ? _canGo_T : _GEN_34; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 124:15 98:18]
  wire  _GEN_39 = 2'h1 == state ? _canIn_T : _GEN_35; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 125:15 98:18]
  wire [38:0] _GEN_41 = 2'h1 == state ? _pnpcOut_T_11 : _GEN_33; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 127:17 98:18]
  wire  canGo = 2'h0 == state ? rvcFinish | rvcNext : _GEN_38; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 100:15 98:18]
  wire  canIn = 2'h0 == state ? rvcFinish | rvcForceLoadNext : _GEN_39; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:15 98:18]
  wire [38:0] pnpcOut = 2'h0 == state ? _pnpcOut_T_5 : _GEN_41; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 103:17 98:18]
  wire  _io_out_bits_brIdx_T_10 = pnpcOut == _pnpcOut_T_9 & _rvcFinish_T_1 | pnpcOut == _pnpcOut_T_7 & isRVC ? 1'h0 : 1'h1
    ; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 185:27]
  assign io_in_ready = ~io_in_valid | _T_11 & canIn | loadNextInstline; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 188:58]
  assign io_out_valid = io_in_valid & canGo; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 187:31]
  assign io_out_bits_instr = {{32'd0}, instr}; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 184:21]
  assign io_out_bits_pc = 2'h0 == state ? io_in_bits_pc : _GEN_40; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 102:15 98:18]
  assign io_out_bits_pnpc = 2'h0 == state ? _pnpcOut_T_5 : _GEN_41; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 103:17 98:18]
  assign io_out_bits_brIdx = {{3'd0}, _io_out_bits_brIdx_T_10}; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 185:21]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 39:22]
      state <= 2'h0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 39:22]
    end else if (~io_flush) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 97:18]
      if (2'h0 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 98:18]
        state <= _GEN_7;
      end else if (2'h1 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 98:18]
        state <= _GEN_7;
      end else begin
        state <= _GEN_36;
      end
    end else begin
      state <= 2'h0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 172:11]
    end
    if (~io_flush) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 97:18]
      if (2'h0 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 98:18]
        specialInstR <= _GEN_10;
      end else if (2'h1 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 98:18]
        specialInstR <= _GEN_10;
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 40:26]
      pcOffsetR <= 3'h0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 40:26]
    end else if (~io_flush) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 97:18]
      if (2'h0 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 98:18]
        pcOffsetR <= _GEN_2;
      end else if (2'h1 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 98:18]
        pcOffsetR <= _GEN_2;
      end else begin
        pcOffsetR <= _GEN_37;
      end
    end
    if (~io_flush) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 97:18]
      if (2'h0 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 98:18]
        specialPCR <= _GEN_8;
      end else if (2'h1 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 98:18]
        specialPCR <= _GEN_8;
      end
    end
    if (~io_flush) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 97:18]
      if (2'h0 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 98:18]
        specialNPCR <= _GEN_9;
      end else if (2'h1 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 98:18]
        specialNPCR <= _GEN_9;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~flushIFU)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at NaiveIBF.scala:59 assert(!flushIFU)\n"); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 59:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  specialInstR = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  pcOffsetR = _RAND_2[2:0];
  _RAND_3 = {2{`RANDOM}};
  specialPCR = _RAND_3[38:0];
  _RAND_4 = {2{`RANDOM}};
  specialNPCR = _RAND_4[38:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (_T_2) begin
      assert(~flushIFU); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 59:9]
    end
  end
endmodule
module Decoder(
  output        io_in_ready, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input         io_in_valid, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input  [63:0] io_in_bits_instr, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input  [38:0] io_in_bits_pc, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input  [38:0] io_in_bits_pnpc, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input  [3:0]  io_in_bits_brIdx, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input         io_out_ready, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_valid, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [63:0] io_out_bits_cf_instr, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [38:0] io_out_bits_cf_pc, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [38:0] io_out_bits_cf_pnpc, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_exceptionVec_1, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_exceptionVec_2, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_0, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_1, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_2, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_3, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_4, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_5, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_6, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_7, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_8, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_9, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_10, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_11, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [3:0]  io_out_bits_cf_brIdx, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_ctrl_src1Type, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_ctrl_src2Type, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [2:0]  io_out_bits_ctrl_fuType, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [6:0]  io_out_bits_ctrl_fuOpType, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [4:0]  io_out_bits_ctrl_rfSrc1, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [4:0]  io_out_bits_ctrl_rfSrc2, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_ctrl_rfWen, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [4:0]  io_out_bits_ctrl_rfDest, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [63:0] io_out_bits_data_imm, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input  [11:0] intrVecIDU
);
  wire [63:0] _decodeList_T = io_in_bits_instr & 64'h707f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_1 = 64'h13 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [63:0] _decodeList_T_2 = io_in_bits_instr & 64'hfc00707f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_3 = 64'h1013 == _decodeList_T_2; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_5 = 64'h2013 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_7 = 64'h3013 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_9 = 64'h4013 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_11 = 64'h5013 == _decodeList_T_2; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_13 = 64'h6013 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_15 = 64'h7013 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_17 = 64'h40005013 == _decodeList_T_2; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [63:0] _decodeList_T_18 = io_in_bits_instr & 64'hfe00707f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_19 = 64'h33 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_21 = 64'h1033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_23 = 64'h2033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_25 = 64'h3033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_27 = 64'h4033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_29 = 64'h5033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_31 = 64'h6033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_33 = 64'h7033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_35 = 64'h40000033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_37 = 64'h40005033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [63:0] _decodeList_T_38 = io_in_bits_instr & 64'h7f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_39 = 64'h17 == _decodeList_T_38; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_41 = 64'h37 == _decodeList_T_38; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_43 = 64'h6f == _decodeList_T_38; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_45 = 64'h67 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_47 = 64'h63 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_49 = 64'h1063 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_51 = 64'h4063 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_53 = 64'h5063 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_55 = 64'h6063 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_57 = 64'h7063 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_59 = 64'h3 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_61 = 64'h1003 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_63 = 64'h2003 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_65 = 64'h4003 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_67 = 64'h5003 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_69 = 64'h23 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_71 = 64'h1023 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_73 = 64'h2023 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_75 = 64'h1b == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_77 = 64'h101b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_79 = 64'h501b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_81 = 64'h4000501b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_83 = 64'h103b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_85 = 64'h503b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_87 = 64'h4000503b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_89 = 64'h3b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_91 = 64'h4000003b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_93 = 64'h6003 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_95 = 64'h3003 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_97 = 64'h3023 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_99 = 64'h6b == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_101 = 64'h2000033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_103 = 64'h2001033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_105 = 64'h2002033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_107 = 64'h2003033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_109 = 64'h2004033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_111 = 64'h2005033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_113 = 64'h2006033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_115 = 64'h2007033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_117 = 64'h200003b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_119 = 64'h200403b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_121 = 64'h200503b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_123 = 64'h200603b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_125 = 64'h200703b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [63:0] _decodeList_T_126 = io_in_bits_instr & 64'hffffffff; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_127 = 64'h73 == _decodeList_T_126; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_129 = 64'h100073 == _decodeList_T_126; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_131 = 64'h30200073 == _decodeList_T_126; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_133 = 64'hf == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_135 = 64'h10500073 == _decodeList_T_126; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [63:0] _decodeList_T_136 = io_in_bits_instr & 64'hf9f0707f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_137 = 64'h1000302f == _decodeList_T_136; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_139 = 64'h1000202f == _decodeList_T_136; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [63:0] _decodeList_T_140 = io_in_bits_instr & 64'hf800707f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_141 = 64'h1800302f == _decodeList_T_140; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_143 = 64'h1800202f == _decodeList_T_140; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [63:0] _decodeList_T_144 = io_in_bits_instr & 64'hf800607f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_145 = 64'h800202f == _decodeList_T_144; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_147 = 64'h202f == _decodeList_T_144; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_149 = 64'h2000202f == _decodeList_T_144; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_151 = 64'h6000202f == _decodeList_T_144; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_153 = 64'h4000202f == _decodeList_T_144; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_155 = 64'h8000202f == _decodeList_T_144; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_157 = 64'ha000202f == _decodeList_T_144; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_159 = 64'hc000202f == _decodeList_T_144; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_161 = 64'he000202f == _decodeList_T_144; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_163 = 64'h1073 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_165 = 64'h2073 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_167 = 64'h3073 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_169 = 64'h5073 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_171 = 64'h6073 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_173 = 64'h7073 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_175 = 64'h100f == _decodeList_T_126; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [2:0] _decodeList_T_177 = _decodeList_T_173 ? 3'h4 : {{2'd0}, _decodeList_T_175}; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_178 = _decodeList_T_171 ? 3'h4 : _decodeList_T_177; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_179 = _decodeList_T_169 ? 3'h4 : _decodeList_T_178; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_180 = _decodeList_T_167 ? 3'h4 : _decodeList_T_179; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_181 = _decodeList_T_165 ? 3'h4 : _decodeList_T_180; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_182 = _decodeList_T_163 ? 3'h4 : _decodeList_T_181; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_183 = _decodeList_T_161 ? 3'h5 : _decodeList_T_182; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_184 = _decodeList_T_159 ? 3'h5 : _decodeList_T_183; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_185 = _decodeList_T_157 ? 3'h5 : _decodeList_T_184; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_186 = _decodeList_T_155 ? 3'h5 : _decodeList_T_185; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_187 = _decodeList_T_153 ? 3'h5 : _decodeList_T_186; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_188 = _decodeList_T_151 ? 3'h5 : _decodeList_T_187; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_189 = _decodeList_T_149 ? 3'h5 : _decodeList_T_188; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_190 = _decodeList_T_147 ? 3'h5 : _decodeList_T_189; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_191 = _decodeList_T_145 ? 3'h5 : _decodeList_T_190; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_192 = _decodeList_T_143 ? 4'hf : {{1'd0}, _decodeList_T_191}; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_193 = _decodeList_T_141 ? 4'hf : _decodeList_T_192; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_194 = _decodeList_T_139 ? 4'h4 : _decodeList_T_193; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_195 = _decodeList_T_137 ? 4'h4 : _decodeList_T_194; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_196 = _decodeList_T_135 ? 4'h4 : _decodeList_T_195; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_197 = _decodeList_T_133 ? 4'h2 : _decodeList_T_196; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_198 = _decodeList_T_131 ? 4'h4 : _decodeList_T_197; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_199 = _decodeList_T_129 ? 4'h4 : _decodeList_T_198; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_200 = _decodeList_T_127 ? 4'h4 : _decodeList_T_199; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_201 = _decodeList_T_125 ? 4'h5 : _decodeList_T_200; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_202 = _decodeList_T_123 ? 4'h5 : _decodeList_T_201; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_203 = _decodeList_T_121 ? 4'h5 : _decodeList_T_202; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_204 = _decodeList_T_119 ? 4'h5 : _decodeList_T_203; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_205 = _decodeList_T_117 ? 4'h5 : _decodeList_T_204; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_206 = _decodeList_T_115 ? 4'h5 : _decodeList_T_205; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_207 = _decodeList_T_113 ? 4'h5 : _decodeList_T_206; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_208 = _decodeList_T_111 ? 4'h5 : _decodeList_T_207; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_209 = _decodeList_T_109 ? 4'h5 : _decodeList_T_208; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_210 = _decodeList_T_107 ? 4'h5 : _decodeList_T_209; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_211 = _decodeList_T_105 ? 4'h5 : _decodeList_T_210; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_212 = _decodeList_T_103 ? 4'h5 : _decodeList_T_211; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_213 = _decodeList_T_101 ? 4'h5 : _decodeList_T_212; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_214 = _decodeList_T_99 ? 4'h4 : _decodeList_T_213; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_215 = _decodeList_T_97 ? 4'h2 : _decodeList_T_214; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_216 = _decodeList_T_95 ? 4'h4 : _decodeList_T_215; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_217 = _decodeList_T_93 ? 4'h4 : _decodeList_T_216; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_218 = _decodeList_T_91 ? 4'h5 : _decodeList_T_217; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_219 = _decodeList_T_89 ? 4'h5 : _decodeList_T_218; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_220 = _decodeList_T_87 ? 4'h5 : _decodeList_T_219; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_221 = _decodeList_T_85 ? 4'h5 : _decodeList_T_220; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_222 = _decodeList_T_83 ? 4'h5 : _decodeList_T_221; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_223 = _decodeList_T_81 ? 4'h4 : _decodeList_T_222; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_224 = _decodeList_T_79 ? 4'h4 : _decodeList_T_223; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_225 = _decodeList_T_77 ? 4'h4 : _decodeList_T_224; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_226 = _decodeList_T_75 ? 4'h4 : _decodeList_T_225; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_227 = _decodeList_T_73 ? 4'h2 : _decodeList_T_226; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_228 = _decodeList_T_71 ? 4'h2 : _decodeList_T_227; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_229 = _decodeList_T_69 ? 4'h2 : _decodeList_T_228; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_230 = _decodeList_T_67 ? 4'h4 : _decodeList_T_229; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_231 = _decodeList_T_65 ? 4'h4 : _decodeList_T_230; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_232 = _decodeList_T_63 ? 4'h4 : _decodeList_T_231; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_233 = _decodeList_T_61 ? 4'h4 : _decodeList_T_232; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_234 = _decodeList_T_59 ? 4'h4 : _decodeList_T_233; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_235 = _decodeList_T_57 ? 4'h1 : _decodeList_T_234; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_236 = _decodeList_T_55 ? 4'h1 : _decodeList_T_235; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_237 = _decodeList_T_53 ? 4'h1 : _decodeList_T_236; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_238 = _decodeList_T_51 ? 4'h1 : _decodeList_T_237; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_239 = _decodeList_T_49 ? 4'h1 : _decodeList_T_238; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_240 = _decodeList_T_47 ? 4'h1 : _decodeList_T_239; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_241 = _decodeList_T_45 ? 4'h4 : _decodeList_T_240; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_242 = _decodeList_T_43 ? 4'h7 : _decodeList_T_241; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_243 = _decodeList_T_41 ? 4'h6 : _decodeList_T_242; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_244 = _decodeList_T_39 ? 4'h6 : _decodeList_T_243; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_245 = _decodeList_T_37 ? 4'h5 : _decodeList_T_244; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_246 = _decodeList_T_35 ? 4'h5 : _decodeList_T_245; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_247 = _decodeList_T_33 ? 4'h5 : _decodeList_T_246; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_248 = _decodeList_T_31 ? 4'h5 : _decodeList_T_247; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_249 = _decodeList_T_29 ? 4'h5 : _decodeList_T_248; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_250 = _decodeList_T_27 ? 4'h5 : _decodeList_T_249; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_251 = _decodeList_T_25 ? 4'h5 : _decodeList_T_250; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_252 = _decodeList_T_23 ? 4'h5 : _decodeList_T_251; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_253 = _decodeList_T_21 ? 4'h5 : _decodeList_T_252; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_254 = _decodeList_T_19 ? 4'h5 : _decodeList_T_253; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_255 = _decodeList_T_17 ? 4'h4 : _decodeList_T_254; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_256 = _decodeList_T_15 ? 4'h4 : _decodeList_T_255; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_257 = _decodeList_T_13 ? 4'h4 : _decodeList_T_256; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_258 = _decodeList_T_11 ? 4'h4 : _decodeList_T_257; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_259 = _decodeList_T_9 ? 4'h4 : _decodeList_T_258; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_260 = _decodeList_T_7 ? 4'h4 : _decodeList_T_259; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_261 = _decodeList_T_5 ? 4'h4 : _decodeList_T_260; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_262 = _decodeList_T_3 ? 4'h4 : _decodeList_T_261; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] decodeList_0 = _decodeList_T_1 ? 4'h4 : _decodeList_T_262; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_263 = _decodeList_T_175 ? 3'h4 : 3'h3; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_264 = _decodeList_T_173 ? 3'h3 : _decodeList_T_263; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_265 = _decodeList_T_171 ? 3'h3 : _decodeList_T_264; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_266 = _decodeList_T_169 ? 3'h3 : _decodeList_T_265; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_267 = _decodeList_T_167 ? 3'h3 : _decodeList_T_266; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_268 = _decodeList_T_165 ? 3'h3 : _decodeList_T_267; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_269 = _decodeList_T_163 ? 3'h3 : _decodeList_T_268; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_270 = _decodeList_T_161 ? 3'h1 : _decodeList_T_269; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_271 = _decodeList_T_159 ? 3'h1 : _decodeList_T_270; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_272 = _decodeList_T_157 ? 3'h1 : _decodeList_T_271; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_273 = _decodeList_T_155 ? 3'h1 : _decodeList_T_272; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_274 = _decodeList_T_153 ? 3'h1 : _decodeList_T_273; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_275 = _decodeList_T_151 ? 3'h1 : _decodeList_T_274; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_276 = _decodeList_T_149 ? 3'h1 : _decodeList_T_275; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_277 = _decodeList_T_147 ? 3'h1 : _decodeList_T_276; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_278 = _decodeList_T_145 ? 3'h1 : _decodeList_T_277; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_279 = _decodeList_T_143 ? 3'h1 : _decodeList_T_278; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_280 = _decodeList_T_141 ? 3'h1 : _decodeList_T_279; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_281 = _decodeList_T_139 ? 3'h1 : _decodeList_T_280; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_282 = _decodeList_T_137 ? 3'h1 : _decodeList_T_281; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_283 = _decodeList_T_135 ? 3'h0 : _decodeList_T_282; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_284 = _decodeList_T_133 ? 3'h4 : _decodeList_T_283; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_285 = _decodeList_T_131 ? 3'h3 : _decodeList_T_284; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_286 = _decodeList_T_129 ? 3'h3 : _decodeList_T_285; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_287 = _decodeList_T_127 ? 3'h3 : _decodeList_T_286; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_288 = _decodeList_T_125 ? 3'h2 : _decodeList_T_287; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_289 = _decodeList_T_123 ? 3'h2 : _decodeList_T_288; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_290 = _decodeList_T_121 ? 3'h2 : _decodeList_T_289; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_291 = _decodeList_T_119 ? 3'h2 : _decodeList_T_290; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_292 = _decodeList_T_117 ? 3'h2 : _decodeList_T_291; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_293 = _decodeList_T_115 ? 3'h2 : _decodeList_T_292; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_294 = _decodeList_T_113 ? 3'h2 : _decodeList_T_293; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_295 = _decodeList_T_111 ? 3'h2 : _decodeList_T_294; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_296 = _decodeList_T_109 ? 3'h2 : _decodeList_T_295; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_297 = _decodeList_T_107 ? 3'h2 : _decodeList_T_296; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_298 = _decodeList_T_105 ? 3'h2 : _decodeList_T_297; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_299 = _decodeList_T_103 ? 3'h2 : _decodeList_T_298; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_300 = _decodeList_T_101 ? 3'h2 : _decodeList_T_299; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_301 = _decodeList_T_99 ? 3'h3 : _decodeList_T_300; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_302 = _decodeList_T_97 ? 3'h1 : _decodeList_T_301; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_303 = _decodeList_T_95 ? 3'h1 : _decodeList_T_302; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_304 = _decodeList_T_93 ? 3'h1 : _decodeList_T_303; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_305 = _decodeList_T_91 ? 3'h0 : _decodeList_T_304; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_306 = _decodeList_T_89 ? 3'h0 : _decodeList_T_305; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_307 = _decodeList_T_87 ? 3'h0 : _decodeList_T_306; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_308 = _decodeList_T_85 ? 3'h0 : _decodeList_T_307; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_309 = _decodeList_T_83 ? 3'h0 : _decodeList_T_308; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_310 = _decodeList_T_81 ? 3'h0 : _decodeList_T_309; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_311 = _decodeList_T_79 ? 3'h0 : _decodeList_T_310; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_312 = _decodeList_T_77 ? 3'h0 : _decodeList_T_311; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_313 = _decodeList_T_75 ? 3'h0 : _decodeList_T_312; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_314 = _decodeList_T_73 ? 3'h1 : _decodeList_T_313; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_315 = _decodeList_T_71 ? 3'h1 : _decodeList_T_314; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_316 = _decodeList_T_69 ? 3'h1 : _decodeList_T_315; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_317 = _decodeList_T_67 ? 3'h1 : _decodeList_T_316; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_318 = _decodeList_T_65 ? 3'h1 : _decodeList_T_317; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_319 = _decodeList_T_63 ? 3'h1 : _decodeList_T_318; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_320 = _decodeList_T_61 ? 3'h1 : _decodeList_T_319; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_321 = _decodeList_T_59 ? 3'h1 : _decodeList_T_320; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_322 = _decodeList_T_57 ? 3'h0 : _decodeList_T_321; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_323 = _decodeList_T_55 ? 3'h0 : _decodeList_T_322; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_324 = _decodeList_T_53 ? 3'h0 : _decodeList_T_323; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_325 = _decodeList_T_51 ? 3'h0 : _decodeList_T_324; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_326 = _decodeList_T_49 ? 3'h0 : _decodeList_T_325; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_327 = _decodeList_T_47 ? 3'h0 : _decodeList_T_326; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_328 = _decodeList_T_45 ? 3'h0 : _decodeList_T_327; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_329 = _decodeList_T_43 ? 3'h0 : _decodeList_T_328; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_330 = _decodeList_T_41 ? 3'h0 : _decodeList_T_329; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_331 = _decodeList_T_39 ? 3'h0 : _decodeList_T_330; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_332 = _decodeList_T_37 ? 3'h0 : _decodeList_T_331; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_333 = _decodeList_T_35 ? 3'h0 : _decodeList_T_332; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_334 = _decodeList_T_33 ? 3'h0 : _decodeList_T_333; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_335 = _decodeList_T_31 ? 3'h0 : _decodeList_T_334; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_336 = _decodeList_T_29 ? 3'h0 : _decodeList_T_335; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_337 = _decodeList_T_27 ? 3'h0 : _decodeList_T_336; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_338 = _decodeList_T_25 ? 3'h0 : _decodeList_T_337; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_339 = _decodeList_T_23 ? 3'h0 : _decodeList_T_338; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_340 = _decodeList_T_21 ? 3'h0 : _decodeList_T_339; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_341 = _decodeList_T_19 ? 3'h0 : _decodeList_T_340; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_342 = _decodeList_T_17 ? 3'h0 : _decodeList_T_341; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_343 = _decodeList_T_15 ? 3'h0 : _decodeList_T_342; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_344 = _decodeList_T_13 ? 3'h0 : _decodeList_T_343; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_345 = _decodeList_T_11 ? 3'h0 : _decodeList_T_344; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_346 = _decodeList_T_9 ? 3'h0 : _decodeList_T_345; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_347 = _decodeList_T_7 ? 3'h0 : _decodeList_T_346; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_348 = _decodeList_T_5 ? 3'h0 : _decodeList_T_347; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_349 = _decodeList_T_3 ? 3'h0 : _decodeList_T_348; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] decodeList_1 = _decodeList_T_1 ? 3'h0 : _decodeList_T_349; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_351 = _decodeList_T_173 ? 3'h7 : {{2'd0}, _decodeList_T_175}; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_352 = _decodeList_T_171 ? 3'h6 : _decodeList_T_351; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_353 = _decodeList_T_169 ? 3'h5 : _decodeList_T_352; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_354 = _decodeList_T_167 ? 3'h3 : _decodeList_T_353; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_355 = _decodeList_T_165 ? 3'h2 : _decodeList_T_354; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_356 = _decodeList_T_163 ? 3'h1 : _decodeList_T_355; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _decodeList_T_357 = _decodeList_T_161 ? 6'h32 : {{3'd0}, _decodeList_T_356}; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _decodeList_T_358 = _decodeList_T_159 ? 6'h31 : _decodeList_T_357; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _decodeList_T_359 = _decodeList_T_157 ? 6'h30 : _decodeList_T_358; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _decodeList_T_360 = _decodeList_T_155 ? 6'h37 : _decodeList_T_359; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _decodeList_T_361 = _decodeList_T_153 ? 6'h26 : _decodeList_T_360; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _decodeList_T_362 = _decodeList_T_151 ? 6'h25 : _decodeList_T_361; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _decodeList_T_363 = _decodeList_T_149 ? 6'h24 : _decodeList_T_362; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_364 = _decodeList_T_147 ? 7'h63 : {{1'd0}, _decodeList_T_363}; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_365 = _decodeList_T_145 ? 7'h22 : _decodeList_T_364; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_366 = _decodeList_T_143 ? 7'h21 : _decodeList_T_365; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_367 = _decodeList_T_141 ? 7'h21 : _decodeList_T_366; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_368 = _decodeList_T_139 ? 7'h20 : _decodeList_T_367; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_369 = _decodeList_T_137 ? 7'h20 : _decodeList_T_368; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_370 = _decodeList_T_135 ? 7'h40 : _decodeList_T_369; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_371 = _decodeList_T_133 ? 7'h0 : _decodeList_T_370; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_372 = _decodeList_T_131 ? 7'h0 : _decodeList_T_371; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_373 = _decodeList_T_129 ? 7'h0 : _decodeList_T_372; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_374 = _decodeList_T_127 ? 7'h0 : _decodeList_T_373; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_375 = _decodeList_T_125 ? 7'hf : _decodeList_T_374; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_376 = _decodeList_T_123 ? 7'he : _decodeList_T_375; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_377 = _decodeList_T_121 ? 7'hd : _decodeList_T_376; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_378 = _decodeList_T_119 ? 7'hc : _decodeList_T_377; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_379 = _decodeList_T_117 ? 7'h8 : _decodeList_T_378; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_380 = _decodeList_T_115 ? 7'h7 : _decodeList_T_379; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_381 = _decodeList_T_113 ? 7'h6 : _decodeList_T_380; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_382 = _decodeList_T_111 ? 7'h5 : _decodeList_T_381; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_383 = _decodeList_T_109 ? 7'h4 : _decodeList_T_382; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_384 = _decodeList_T_107 ? 7'h3 : _decodeList_T_383; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_385 = _decodeList_T_105 ? 7'h2 : _decodeList_T_384; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_386 = _decodeList_T_103 ? 7'h1 : _decodeList_T_385; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_387 = _decodeList_T_101 ? 7'h0 : _decodeList_T_386; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_388 = _decodeList_T_99 ? 7'h2 : _decodeList_T_387; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_389 = _decodeList_T_97 ? 7'hb : _decodeList_T_388; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_390 = _decodeList_T_95 ? 7'h3 : _decodeList_T_389; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_391 = _decodeList_T_93 ? 7'h6 : _decodeList_T_390; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_392 = _decodeList_T_91 ? 7'h28 : _decodeList_T_391; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_393 = _decodeList_T_89 ? 7'h60 : _decodeList_T_392; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_394 = _decodeList_T_87 ? 7'h2d : _decodeList_T_393; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_395 = _decodeList_T_85 ? 7'h25 : _decodeList_T_394; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_396 = _decodeList_T_83 ? 7'h21 : _decodeList_T_395; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_397 = _decodeList_T_81 ? 7'h2d : _decodeList_T_396; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_398 = _decodeList_T_79 ? 7'h25 : _decodeList_T_397; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_399 = _decodeList_T_77 ? 7'h21 : _decodeList_T_398; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_400 = _decodeList_T_75 ? 7'h60 : _decodeList_T_399; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_401 = _decodeList_T_73 ? 7'ha : _decodeList_T_400; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_402 = _decodeList_T_71 ? 7'h9 : _decodeList_T_401; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_403 = _decodeList_T_69 ? 7'h8 : _decodeList_T_402; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_404 = _decodeList_T_67 ? 7'h5 : _decodeList_T_403; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_405 = _decodeList_T_65 ? 7'h4 : _decodeList_T_404; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_406 = _decodeList_T_63 ? 7'h2 : _decodeList_T_405; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_407 = _decodeList_T_61 ? 7'h1 : _decodeList_T_406; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_408 = _decodeList_T_59 ? 7'h0 : _decodeList_T_407; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_409 = _decodeList_T_57 ? 7'h17 : _decodeList_T_408; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_410 = _decodeList_T_55 ? 7'h16 : _decodeList_T_409; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_411 = _decodeList_T_53 ? 7'h15 : _decodeList_T_410; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_412 = _decodeList_T_51 ? 7'h14 : _decodeList_T_411; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_413 = _decodeList_T_49 ? 7'h11 : _decodeList_T_412; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_414 = _decodeList_T_47 ? 7'h10 : _decodeList_T_413; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_415 = _decodeList_T_45 ? 7'h5a : _decodeList_T_414; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_416 = _decodeList_T_43 ? 7'h58 : _decodeList_T_415; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_417 = _decodeList_T_41 ? 7'h40 : _decodeList_T_416; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_418 = _decodeList_T_39 ? 7'h40 : _decodeList_T_417; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_419 = _decodeList_T_37 ? 7'hd : _decodeList_T_418; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_420 = _decodeList_T_35 ? 7'hb : _decodeList_T_419; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_421 = _decodeList_T_33 ? 7'h7 : _decodeList_T_420; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_422 = _decodeList_T_31 ? 7'h6 : _decodeList_T_421; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_423 = _decodeList_T_29 ? 7'h5 : _decodeList_T_422; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_424 = _decodeList_T_27 ? 7'h4 : _decodeList_T_423; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_425 = _decodeList_T_25 ? 7'h3 : _decodeList_T_424; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_426 = _decodeList_T_23 ? 7'h2 : _decodeList_T_425; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_427 = _decodeList_T_21 ? 7'h1 : _decodeList_T_426; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_428 = _decodeList_T_19 ? 7'h40 : _decodeList_T_427; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_429 = _decodeList_T_17 ? 7'hd : _decodeList_T_428; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_430 = _decodeList_T_15 ? 7'h7 : _decodeList_T_429; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_431 = _decodeList_T_13 ? 7'h6 : _decodeList_T_430; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_432 = _decodeList_T_11 ? 7'h5 : _decodeList_T_431; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_433 = _decodeList_T_9 ? 7'h4 : _decodeList_T_432; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_434 = _decodeList_T_7 ? 7'h3 : _decodeList_T_433; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_435 = _decodeList_T_5 ? 7'h2 : _decodeList_T_434; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_436 = _decodeList_T_3 ? 7'h1 : _decodeList_T_435; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] decodeList_2 = _decodeList_T_1 ? 7'h40 : _decodeList_T_436; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  hasIntr = |intrVecIDU; // @[src/main/scala/nutcore/frontend/IDU.scala 172:22]
  wire [3:0] instrType = hasIntr | io_out_bits_cf_exceptionVec_1 ? 4'h0 : decodeList_0; // @[src/main/scala/nutcore/frontend/IDU.scala 38:75]
  wire [2:0] fuType = hasIntr | io_out_bits_cf_exceptionVec_1 ? 3'h3 : decodeList_1; // @[src/main/scala/nutcore/frontend/IDU.scala 38:75]
  wire [6:0] fuOpType = hasIntr | io_out_bits_cf_exceptionVec_1 ? 7'h0 : decodeList_2; // @[src/main/scala/nutcore/frontend/IDU.scala 38:75]
  wire  _src1Type_T = 4'h4 == instrType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _src1Type_T_2 = 4'h2 == instrType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _src1Type_T_3 = 4'hf == instrType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _src1Type_T_4 = 4'h1 == instrType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _src1Type_T_5 = 4'h6 == instrType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _src1Type_T_6 = 4'h7 == instrType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _src1Type_T_7 = 4'h0 == instrType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  src1Type = _src1Type_T_5 | _src1Type_T_6 | _src1Type_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  src2Type = _src1Type_T | _src1Type_T_5 | _src1Type_T_6 | _src1Type_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] rs = io_in_bits_instr[19:15]; // @[src/main/scala/nutcore/frontend/IDU.scala 62:28]
  wire [4:0] rt = io_in_bits_instr[24:20]; // @[src/main/scala/nutcore/frontend/IDU.scala 62:43]
  wire [4:0] rd = io_in_bits_instr[11:7]; // @[src/main/scala/nutcore/frontend/IDU.scala 62:58]
  wire  imm_signBit = io_in_bits_instr[31]; // @[src/main/scala/utils/BitUtils.scala 39:20]
  wire [51:0] _imm_T_2 = imm_signBit ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/utils/BitUtils.scala 40:46]
  wire [63:0] _imm_T_3 = {_imm_T_2,io_in_bits_instr[31:20]}; // @[src/main/scala/utils/BitUtils.scala 40:41]
  wire [11:0] _imm_T_6 = {io_in_bits_instr[31:25],rd}; // @[src/main/scala/nutcore/frontend/IDU.scala 102:27]
  wire  imm_signBit_1 = _imm_T_6[11]; // @[src/main/scala/utils/BitUtils.scala 39:20]
  wire [51:0] _imm_T_8 = imm_signBit_1 ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/utils/BitUtils.scala 40:46]
  wire [63:0] _imm_T_9 = {_imm_T_8,io_in_bits_instr[31:25],rd}; // @[src/main/scala/utils/BitUtils.scala 40:41]
  wire [12:0] _imm_T_20 = {io_in_bits_instr[31],io_in_bits_instr[7],io_in_bits_instr[30:25],io_in_bits_instr[11:8],1'h0}
    ; // @[src/main/scala/nutcore/frontend/IDU.scala 104:27]
  wire  imm_signBit_3 = _imm_T_20[12]; // @[src/main/scala/utils/BitUtils.scala 39:20]
  wire [50:0] _imm_T_22 = imm_signBit_3 ? 51'h7ffffffffffff : 51'h0; // @[src/main/scala/utils/BitUtils.scala 40:46]
  wire [63:0] _imm_T_23 = {_imm_T_22,io_in_bits_instr[31],io_in_bits_instr[7],io_in_bits_instr[30:25],io_in_bits_instr[
    11:8],1'h0}; // @[src/main/scala/utils/BitUtils.scala 40:41]
  wire [31:0] _imm_T_25 = {io_in_bits_instr[31:12],12'h0}; // @[src/main/scala/nutcore/frontend/IDU.scala 105:27]
  wire  imm_signBit_4 = _imm_T_25[31]; // @[src/main/scala/utils/BitUtils.scala 39:20]
  wire [31:0] _imm_T_27 = imm_signBit_4 ? 32'hffffffff : 32'h0; // @[src/main/scala/utils/BitUtils.scala 40:46]
  wire [63:0] _imm_T_28 = {_imm_T_27,io_in_bits_instr[31:12],12'h0}; // @[src/main/scala/utils/BitUtils.scala 40:41]
  wire [20:0] _imm_T_33 = {io_in_bits_instr[31],io_in_bits_instr[19:12],io_in_bits_instr[20],io_in_bits_instr[30:21],1'h0
    }; // @[src/main/scala/nutcore/frontend/IDU.scala 106:27]
  wire  imm_signBit_5 = _imm_T_33[20]; // @[src/main/scala/utils/BitUtils.scala 39:20]
  wire [42:0] _imm_T_35 = imm_signBit_5 ? 43'h7ffffffffff : 43'h0; // @[src/main/scala/utils/BitUtils.scala 40:46]
  wire [63:0] _imm_T_36 = {_imm_T_35,io_in_bits_instr[31],io_in_bits_instr[19:12],io_in_bits_instr[20],io_in_bits_instr[
    30:21],1'h0}; // @[src/main/scala/utils/BitUtils.scala 40:41]
  wire [63:0] _imm_T_43 = _src1Type_T ? _imm_T_3 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_44 = _src1Type_T_2 ? _imm_T_9 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_45 = _src1Type_T_3 ? _imm_T_9 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_46 = _src1Type_T_4 ? _imm_T_23 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_47 = _src1Type_T_5 ? _imm_T_28 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_48 = _src1Type_T_6 ? _imm_T_36 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_49 = _imm_T_43 | _imm_T_44; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_50 = _imm_T_49 | _imm_T_45; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_51 = _imm_T_50 | _imm_T_46; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_52 = _imm_T_51 | _imm_T_47; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _T_203 = rd == 5'h1 | rd == 5'h5; // @[src/main/scala/nutcore/frontend/IDU.scala 133:42]
  wire [6:0] _GEN_0 = _T_203 & fuOpType == 7'h58 ? 7'h5c : fuOpType; // @[src/main/scala/nutcore/frontend/IDU.scala 134:{57,85} 47:29]
  wire  _T_209 = rs == 5'h1 | rs == 5'h5; // @[src/main/scala/nutcore/frontend/IDU.scala 133:42]
  wire [6:0] _GEN_1 = _T_209 ? 7'h5e : _GEN_0; // @[src/main/scala/nutcore/frontend/IDU.scala 136:{29,57}]
  wire [6:0] _GEN_2 = _T_203 ? 7'h5c : _GEN_1; // @[src/main/scala/nutcore/frontend/IDU.scala 137:{29,57}]
  wire [6:0] _GEN_3 = fuOpType == 7'h5a ? _GEN_2 : _GEN_0; // @[src/main/scala/nutcore/frontend/IDU.scala 135:40]
  wire  _io_in_ready_T_1 = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _io_in_ready_T_2 = ~hasIntr; // @[src/main/scala/nutcore/frontend/IDU.scala 162:49]
  assign io_in_ready = ~io_in_valid | _io_in_ready_T_1 & ~hasIntr; // @[src/main/scala/nutcore/frontend/IDU.scala 162:31]
  assign io_out_valid = io_in_valid; // @[src/main/scala/nutcore/frontend/IDU.scala 161:16]
  assign io_out_bits_cf_instr = io_in_bits_instr; // @[src/main/scala/nutcore/frontend/IDU.scala 163:18]
  assign io_out_bits_cf_pc = io_in_bits_pc; // @[src/main/scala/nutcore/frontend/IDU.scala 163:18]
  assign io_out_bits_cf_pnpc = io_in_bits_pnpc; // @[src/main/scala/nutcore/frontend/IDU.scala 163:18]
  assign io_out_bits_cf_exceptionVec_1 = |io_in_bits_pc[38:32]; // @[src/main/scala/nutcore/frontend/IDU.scala 190:94]
  assign io_out_bits_cf_exceptionVec_2 = instrType == 4'h0 & _io_in_ready_T_2 & io_in_valid; // @[src/main/scala/nutcore/frontend/IDU.scala 178:83]
  assign io_out_bits_cf_intrVec_0 = intrVecIDU[0]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_1 = intrVecIDU[1]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_2 = intrVecIDU[2]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_3 = intrVecIDU[3]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_4 = intrVecIDU[4]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_5 = intrVecIDU[5]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_6 = intrVecIDU[6]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_7 = intrVecIDU[7]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_8 = intrVecIDU[8]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_9 = intrVecIDU[9]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_10 = intrVecIDU[10]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_11 = intrVecIDU[11]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_brIdx = io_in_bits_brIdx; // @[src/main/scala/nutcore/frontend/IDU.scala 163:18]
  assign io_out_bits_ctrl_src1Type = io_in_bits_instr[6:0] == 7'h37 ? 1'h0 : src1Type; // @[src/main/scala/nutcore/frontend/IDU.scala 141:35]
  assign io_out_bits_ctrl_src2Type = _src1Type_T | _src1Type_T_5 | _src1Type_T_6 | _src1Type_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_out_bits_ctrl_fuType = hasIntr | io_out_bits_cf_exceptionVec_1 ? 3'h3 : decodeList_1; // @[src/main/scala/nutcore/frontend/IDU.scala 38:75]
  assign io_out_bits_ctrl_fuOpType = fuType == 3'h0 ? _GEN_3 : fuOpType; // @[src/main/scala/nutcore/frontend/IDU.scala 132:32 47:29]
  assign io_out_bits_ctrl_rfSrc1 = src1Type ? 5'h0 : rs; // @[src/main/scala/nutcore/frontend/IDU.scala 94:33]
  assign io_out_bits_ctrl_rfSrc2 = ~src2Type ? rt : 5'h0; // @[src/main/scala/nutcore/frontend/IDU.scala 95:33]
  assign io_out_bits_ctrl_rfWen = instrType[2]; // @[src/main/scala/nutcore/Decode.scala 33:50]
  assign io_out_bits_ctrl_rfDest = instrType[2] ? rd : 5'h0; // @[src/main/scala/nutcore/frontend/IDU.scala 97:33]
  assign io_out_bits_data_imm = _imm_T_52 | _imm_T_48; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
endmodule
module Decoder_1(
  output        io_out_bits_cf_intrVec_0, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_1, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_2, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_3, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_4, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_5, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_6, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_7, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_8, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_9, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_10, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_11, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input  [11:0] intrVecIDU
);
  assign io_out_bits_cf_intrVec_0 = intrVecIDU[0]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_1 = intrVecIDU[1]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_2 = intrVecIDU[2]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_3 = intrVecIDU[3]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_4 = intrVecIDU[4]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_5 = intrVecIDU[5]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_6 = intrVecIDU[6]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_7 = intrVecIDU[7]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_8 = intrVecIDU[8]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_9 = intrVecIDU[9]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_10 = intrVecIDU[10]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
  assign io_out_bits_cf_intrVec_11 = intrVecIDU[11]; // @[src/main/scala/nutcore/frontend/IDU.scala 171:38]
endmodule
module IDU(
  output        io_in_0_ready, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  input         io_in_0_valid, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  input  [63:0] io_in_0_bits_instr, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  input  [38:0] io_in_0_bits_pc, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  input  [38:0] io_in_0_bits_pnpc, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  input  [3:0]  io_in_0_bits_brIdx, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  input         io_out_0_ready, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  output        io_out_0_valid, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  output [63:0] io_out_0_bits_cf_instr, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  output [38:0] io_out_0_bits_cf_pc, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  output [38:0] io_out_0_bits_cf_pnpc, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  output        io_out_0_bits_cf_exceptionVec_1, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  output        io_out_0_bits_cf_exceptionVec_2, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  output        io_out_0_bits_cf_intrVec_0, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  output        io_out_0_bits_cf_intrVec_1, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  output        io_out_0_bits_cf_intrVec_2, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  output        io_out_0_bits_cf_intrVec_3, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  output        io_out_0_bits_cf_intrVec_4, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  output        io_out_0_bits_cf_intrVec_5, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  output        io_out_0_bits_cf_intrVec_6, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  output        io_out_0_bits_cf_intrVec_7, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  output        io_out_0_bits_cf_intrVec_8, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  output        io_out_0_bits_cf_intrVec_9, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  output        io_out_0_bits_cf_intrVec_10, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  output        io_out_0_bits_cf_intrVec_11, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  output [3:0]  io_out_0_bits_cf_brIdx, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  output        io_out_0_bits_ctrl_src1Type, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  output        io_out_0_bits_ctrl_src2Type, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  output [2:0]  io_out_0_bits_ctrl_fuType, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  output [6:0]  io_out_0_bits_ctrl_fuOpType, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  output [4:0]  io_out_0_bits_ctrl_rfSrc1, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  output [4:0]  io_out_0_bits_ctrl_rfSrc2, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  output        io_out_0_bits_ctrl_rfWen, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  output [4:0]  io_out_0_bits_ctrl_rfDest, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  output [63:0] io_out_0_bits_data_imm, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  output        io_out_1_bits_cf_intrVec_0, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  output        io_out_1_bits_cf_intrVec_1, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  output        io_out_1_bits_cf_intrVec_2, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  output        io_out_1_bits_cf_intrVec_3, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  output        io_out_1_bits_cf_intrVec_4, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  output        io_out_1_bits_cf_intrVec_5, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  output        io_out_1_bits_cf_intrVec_6, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  output        io_out_1_bits_cf_intrVec_7, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  output        io_out_1_bits_cf_intrVec_8, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  output        io_out_1_bits_cf_intrVec_9, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  output        io_out_1_bits_cf_intrVec_10, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  output        io_out_1_bits_cf_intrVec_11, // @[src/main/scala/nutcore/frontend/IDU.scala 202:14]
  input  [11:0] intrVec
);
  wire  decoder1_io_in_ready; // @[src/main/scala/nutcore/frontend/IDU.scala 206:25]
  wire  decoder1_io_in_valid; // @[src/main/scala/nutcore/frontend/IDU.scala 206:25]
  wire [63:0] decoder1_io_in_bits_instr; // @[src/main/scala/nutcore/frontend/IDU.scala 206:25]
  wire [38:0] decoder1_io_in_bits_pc; // @[src/main/scala/nutcore/frontend/IDU.scala 206:25]
  wire [38:0] decoder1_io_in_bits_pnpc; // @[src/main/scala/nutcore/frontend/IDU.scala 206:25]
  wire [3:0] decoder1_io_in_bits_brIdx; // @[src/main/scala/nutcore/frontend/IDU.scala 206:25]
  wire  decoder1_io_out_ready; // @[src/main/scala/nutcore/frontend/IDU.scala 206:25]
  wire  decoder1_io_out_valid; // @[src/main/scala/nutcore/frontend/IDU.scala 206:25]
  wire [63:0] decoder1_io_out_bits_cf_instr; // @[src/main/scala/nutcore/frontend/IDU.scala 206:25]
  wire [38:0] decoder1_io_out_bits_cf_pc; // @[src/main/scala/nutcore/frontend/IDU.scala 206:25]
  wire [38:0] decoder1_io_out_bits_cf_pnpc; // @[src/main/scala/nutcore/frontend/IDU.scala 206:25]
  wire  decoder1_io_out_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/frontend/IDU.scala 206:25]
  wire  decoder1_io_out_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/frontend/IDU.scala 206:25]
  wire  decoder1_io_out_bits_cf_intrVec_0; // @[src/main/scala/nutcore/frontend/IDU.scala 206:25]
  wire  decoder1_io_out_bits_cf_intrVec_1; // @[src/main/scala/nutcore/frontend/IDU.scala 206:25]
  wire  decoder1_io_out_bits_cf_intrVec_2; // @[src/main/scala/nutcore/frontend/IDU.scala 206:25]
  wire  decoder1_io_out_bits_cf_intrVec_3; // @[src/main/scala/nutcore/frontend/IDU.scala 206:25]
  wire  decoder1_io_out_bits_cf_intrVec_4; // @[src/main/scala/nutcore/frontend/IDU.scala 206:25]
  wire  decoder1_io_out_bits_cf_intrVec_5; // @[src/main/scala/nutcore/frontend/IDU.scala 206:25]
  wire  decoder1_io_out_bits_cf_intrVec_6; // @[src/main/scala/nutcore/frontend/IDU.scala 206:25]
  wire  decoder1_io_out_bits_cf_intrVec_7; // @[src/main/scala/nutcore/frontend/IDU.scala 206:25]
  wire  decoder1_io_out_bits_cf_intrVec_8; // @[src/main/scala/nutcore/frontend/IDU.scala 206:25]
  wire  decoder1_io_out_bits_cf_intrVec_9; // @[src/main/scala/nutcore/frontend/IDU.scala 206:25]
  wire  decoder1_io_out_bits_cf_intrVec_10; // @[src/main/scala/nutcore/frontend/IDU.scala 206:25]
  wire  decoder1_io_out_bits_cf_intrVec_11; // @[src/main/scala/nutcore/frontend/IDU.scala 206:25]
  wire [3:0] decoder1_io_out_bits_cf_brIdx; // @[src/main/scala/nutcore/frontend/IDU.scala 206:25]
  wire  decoder1_io_out_bits_ctrl_src1Type; // @[src/main/scala/nutcore/frontend/IDU.scala 206:25]
  wire  decoder1_io_out_bits_ctrl_src2Type; // @[src/main/scala/nutcore/frontend/IDU.scala 206:25]
  wire [2:0] decoder1_io_out_bits_ctrl_fuType; // @[src/main/scala/nutcore/frontend/IDU.scala 206:25]
  wire [6:0] decoder1_io_out_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/frontend/IDU.scala 206:25]
  wire [4:0] decoder1_io_out_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/frontend/IDU.scala 206:25]
  wire [4:0] decoder1_io_out_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/frontend/IDU.scala 206:25]
  wire  decoder1_io_out_bits_ctrl_rfWen; // @[src/main/scala/nutcore/frontend/IDU.scala 206:25]
  wire [4:0] decoder1_io_out_bits_ctrl_rfDest; // @[src/main/scala/nutcore/frontend/IDU.scala 206:25]
  wire [63:0] decoder1_io_out_bits_data_imm; // @[src/main/scala/nutcore/frontend/IDU.scala 206:25]
  wire [11:0] decoder1_intrVecIDU; // @[src/main/scala/nutcore/frontend/IDU.scala 206:25]
  wire  decoder2_io_out_bits_cf_intrVec_0; // @[src/main/scala/nutcore/frontend/IDU.scala 207:25]
  wire  decoder2_io_out_bits_cf_intrVec_1; // @[src/main/scala/nutcore/frontend/IDU.scala 207:25]
  wire  decoder2_io_out_bits_cf_intrVec_2; // @[src/main/scala/nutcore/frontend/IDU.scala 207:25]
  wire  decoder2_io_out_bits_cf_intrVec_3; // @[src/main/scala/nutcore/frontend/IDU.scala 207:25]
  wire  decoder2_io_out_bits_cf_intrVec_4; // @[src/main/scala/nutcore/frontend/IDU.scala 207:25]
  wire  decoder2_io_out_bits_cf_intrVec_5; // @[src/main/scala/nutcore/frontend/IDU.scala 207:25]
  wire  decoder2_io_out_bits_cf_intrVec_6; // @[src/main/scala/nutcore/frontend/IDU.scala 207:25]
  wire  decoder2_io_out_bits_cf_intrVec_7; // @[src/main/scala/nutcore/frontend/IDU.scala 207:25]
  wire  decoder2_io_out_bits_cf_intrVec_8; // @[src/main/scala/nutcore/frontend/IDU.scala 207:25]
  wire  decoder2_io_out_bits_cf_intrVec_9; // @[src/main/scala/nutcore/frontend/IDU.scala 207:25]
  wire  decoder2_io_out_bits_cf_intrVec_10; // @[src/main/scala/nutcore/frontend/IDU.scala 207:25]
  wire  decoder2_io_out_bits_cf_intrVec_11; // @[src/main/scala/nutcore/frontend/IDU.scala 207:25]
  wire [11:0] decoder2_intrVecIDU; // @[src/main/scala/nutcore/frontend/IDU.scala 207:25]
  Decoder decoder1 ( // @[src/main/scala/nutcore/frontend/IDU.scala 206:25]
    .io_in_ready(decoder1_io_in_ready),
    .io_in_valid(decoder1_io_in_valid),
    .io_in_bits_instr(decoder1_io_in_bits_instr),
    .io_in_bits_pc(decoder1_io_in_bits_pc),
    .io_in_bits_pnpc(decoder1_io_in_bits_pnpc),
    .io_in_bits_brIdx(decoder1_io_in_bits_brIdx),
    .io_out_ready(decoder1_io_out_ready),
    .io_out_valid(decoder1_io_out_valid),
    .io_out_bits_cf_instr(decoder1_io_out_bits_cf_instr),
    .io_out_bits_cf_pc(decoder1_io_out_bits_cf_pc),
    .io_out_bits_cf_pnpc(decoder1_io_out_bits_cf_pnpc),
    .io_out_bits_cf_exceptionVec_1(decoder1_io_out_bits_cf_exceptionVec_1),
    .io_out_bits_cf_exceptionVec_2(decoder1_io_out_bits_cf_exceptionVec_2),
    .io_out_bits_cf_intrVec_0(decoder1_io_out_bits_cf_intrVec_0),
    .io_out_bits_cf_intrVec_1(decoder1_io_out_bits_cf_intrVec_1),
    .io_out_bits_cf_intrVec_2(decoder1_io_out_bits_cf_intrVec_2),
    .io_out_bits_cf_intrVec_3(decoder1_io_out_bits_cf_intrVec_3),
    .io_out_bits_cf_intrVec_4(decoder1_io_out_bits_cf_intrVec_4),
    .io_out_bits_cf_intrVec_5(decoder1_io_out_bits_cf_intrVec_5),
    .io_out_bits_cf_intrVec_6(decoder1_io_out_bits_cf_intrVec_6),
    .io_out_bits_cf_intrVec_7(decoder1_io_out_bits_cf_intrVec_7),
    .io_out_bits_cf_intrVec_8(decoder1_io_out_bits_cf_intrVec_8),
    .io_out_bits_cf_intrVec_9(decoder1_io_out_bits_cf_intrVec_9),
    .io_out_bits_cf_intrVec_10(decoder1_io_out_bits_cf_intrVec_10),
    .io_out_bits_cf_intrVec_11(decoder1_io_out_bits_cf_intrVec_11),
    .io_out_bits_cf_brIdx(decoder1_io_out_bits_cf_brIdx),
    .io_out_bits_ctrl_src1Type(decoder1_io_out_bits_ctrl_src1Type),
    .io_out_bits_ctrl_src2Type(decoder1_io_out_bits_ctrl_src2Type),
    .io_out_bits_ctrl_fuType(decoder1_io_out_bits_ctrl_fuType),
    .io_out_bits_ctrl_fuOpType(decoder1_io_out_bits_ctrl_fuOpType),
    .io_out_bits_ctrl_rfSrc1(decoder1_io_out_bits_ctrl_rfSrc1),
    .io_out_bits_ctrl_rfSrc2(decoder1_io_out_bits_ctrl_rfSrc2),
    .io_out_bits_ctrl_rfWen(decoder1_io_out_bits_ctrl_rfWen),
    .io_out_bits_ctrl_rfDest(decoder1_io_out_bits_ctrl_rfDest),
    .io_out_bits_data_imm(decoder1_io_out_bits_data_imm),
    .intrVecIDU(decoder1_intrVecIDU)
  );
  Decoder_1 decoder2 ( // @[src/main/scala/nutcore/frontend/IDU.scala 207:25]
    .io_out_bits_cf_intrVec_0(decoder2_io_out_bits_cf_intrVec_0),
    .io_out_bits_cf_intrVec_1(decoder2_io_out_bits_cf_intrVec_1),
    .io_out_bits_cf_intrVec_2(decoder2_io_out_bits_cf_intrVec_2),
    .io_out_bits_cf_intrVec_3(decoder2_io_out_bits_cf_intrVec_3),
    .io_out_bits_cf_intrVec_4(decoder2_io_out_bits_cf_intrVec_4),
    .io_out_bits_cf_intrVec_5(decoder2_io_out_bits_cf_intrVec_5),
    .io_out_bits_cf_intrVec_6(decoder2_io_out_bits_cf_intrVec_6),
    .io_out_bits_cf_intrVec_7(decoder2_io_out_bits_cf_intrVec_7),
    .io_out_bits_cf_intrVec_8(decoder2_io_out_bits_cf_intrVec_8),
    .io_out_bits_cf_intrVec_9(decoder2_io_out_bits_cf_intrVec_9),
    .io_out_bits_cf_intrVec_10(decoder2_io_out_bits_cf_intrVec_10),
    .io_out_bits_cf_intrVec_11(decoder2_io_out_bits_cf_intrVec_11),
    .intrVecIDU(decoder2_intrVecIDU)
  );
  assign io_in_0_ready = decoder1_io_in_ready; // @[src/main/scala/nutcore/frontend/IDU.scala 208:12]
  assign io_out_0_valid = decoder1_io_out_valid; // @[src/main/scala/nutcore/frontend/IDU.scala 210:13]
  assign io_out_0_bits_cf_instr = decoder1_io_out_bits_cf_instr; // @[src/main/scala/nutcore/frontend/IDU.scala 210:13]
  assign io_out_0_bits_cf_pc = decoder1_io_out_bits_cf_pc; // @[src/main/scala/nutcore/frontend/IDU.scala 210:13]
  assign io_out_0_bits_cf_pnpc = decoder1_io_out_bits_cf_pnpc; // @[src/main/scala/nutcore/frontend/IDU.scala 210:13]
  assign io_out_0_bits_cf_exceptionVec_1 = decoder1_io_out_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/frontend/IDU.scala 210:13]
  assign io_out_0_bits_cf_exceptionVec_2 = decoder1_io_out_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/frontend/IDU.scala 210:13]
  assign io_out_0_bits_cf_intrVec_0 = decoder1_io_out_bits_cf_intrVec_0; // @[src/main/scala/nutcore/frontend/IDU.scala 210:13]
  assign io_out_0_bits_cf_intrVec_1 = decoder1_io_out_bits_cf_intrVec_1; // @[src/main/scala/nutcore/frontend/IDU.scala 210:13]
  assign io_out_0_bits_cf_intrVec_2 = decoder1_io_out_bits_cf_intrVec_2; // @[src/main/scala/nutcore/frontend/IDU.scala 210:13]
  assign io_out_0_bits_cf_intrVec_3 = decoder1_io_out_bits_cf_intrVec_3; // @[src/main/scala/nutcore/frontend/IDU.scala 210:13]
  assign io_out_0_bits_cf_intrVec_4 = decoder1_io_out_bits_cf_intrVec_4; // @[src/main/scala/nutcore/frontend/IDU.scala 210:13]
  assign io_out_0_bits_cf_intrVec_5 = decoder1_io_out_bits_cf_intrVec_5; // @[src/main/scala/nutcore/frontend/IDU.scala 210:13]
  assign io_out_0_bits_cf_intrVec_6 = decoder1_io_out_bits_cf_intrVec_6; // @[src/main/scala/nutcore/frontend/IDU.scala 210:13]
  assign io_out_0_bits_cf_intrVec_7 = decoder1_io_out_bits_cf_intrVec_7; // @[src/main/scala/nutcore/frontend/IDU.scala 210:13]
  assign io_out_0_bits_cf_intrVec_8 = decoder1_io_out_bits_cf_intrVec_8; // @[src/main/scala/nutcore/frontend/IDU.scala 210:13]
  assign io_out_0_bits_cf_intrVec_9 = decoder1_io_out_bits_cf_intrVec_9; // @[src/main/scala/nutcore/frontend/IDU.scala 210:13]
  assign io_out_0_bits_cf_intrVec_10 = decoder1_io_out_bits_cf_intrVec_10; // @[src/main/scala/nutcore/frontend/IDU.scala 210:13]
  assign io_out_0_bits_cf_intrVec_11 = decoder1_io_out_bits_cf_intrVec_11; // @[src/main/scala/nutcore/frontend/IDU.scala 210:13]
  assign io_out_0_bits_cf_brIdx = decoder1_io_out_bits_cf_brIdx; // @[src/main/scala/nutcore/frontend/IDU.scala 210:13]
  assign io_out_0_bits_ctrl_src1Type = decoder1_io_out_bits_ctrl_src1Type; // @[src/main/scala/nutcore/frontend/IDU.scala 210:13]
  assign io_out_0_bits_ctrl_src2Type = decoder1_io_out_bits_ctrl_src2Type; // @[src/main/scala/nutcore/frontend/IDU.scala 210:13]
  assign io_out_0_bits_ctrl_fuType = decoder1_io_out_bits_ctrl_fuType; // @[src/main/scala/nutcore/frontend/IDU.scala 210:13]
  assign io_out_0_bits_ctrl_fuOpType = decoder1_io_out_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/frontend/IDU.scala 210:13]
  assign io_out_0_bits_ctrl_rfSrc1 = decoder1_io_out_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/frontend/IDU.scala 210:13]
  assign io_out_0_bits_ctrl_rfSrc2 = decoder1_io_out_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/frontend/IDU.scala 210:13]
  assign io_out_0_bits_ctrl_rfWen = decoder1_io_out_bits_ctrl_rfWen; // @[src/main/scala/nutcore/frontend/IDU.scala 210:13]
  assign io_out_0_bits_ctrl_rfDest = decoder1_io_out_bits_ctrl_rfDest; // @[src/main/scala/nutcore/frontend/IDU.scala 210:13]
  assign io_out_0_bits_data_imm = decoder1_io_out_bits_data_imm; // @[src/main/scala/nutcore/frontend/IDU.scala 210:13]
  assign io_out_1_bits_cf_intrVec_0 = decoder2_io_out_bits_cf_intrVec_0; // @[src/main/scala/nutcore/frontend/IDU.scala 211:13]
  assign io_out_1_bits_cf_intrVec_1 = decoder2_io_out_bits_cf_intrVec_1; // @[src/main/scala/nutcore/frontend/IDU.scala 211:13]
  assign io_out_1_bits_cf_intrVec_2 = decoder2_io_out_bits_cf_intrVec_2; // @[src/main/scala/nutcore/frontend/IDU.scala 211:13]
  assign io_out_1_bits_cf_intrVec_3 = decoder2_io_out_bits_cf_intrVec_3; // @[src/main/scala/nutcore/frontend/IDU.scala 211:13]
  assign io_out_1_bits_cf_intrVec_4 = decoder2_io_out_bits_cf_intrVec_4; // @[src/main/scala/nutcore/frontend/IDU.scala 211:13]
  assign io_out_1_bits_cf_intrVec_5 = decoder2_io_out_bits_cf_intrVec_5; // @[src/main/scala/nutcore/frontend/IDU.scala 211:13]
  assign io_out_1_bits_cf_intrVec_6 = decoder2_io_out_bits_cf_intrVec_6; // @[src/main/scala/nutcore/frontend/IDU.scala 211:13]
  assign io_out_1_bits_cf_intrVec_7 = decoder2_io_out_bits_cf_intrVec_7; // @[src/main/scala/nutcore/frontend/IDU.scala 211:13]
  assign io_out_1_bits_cf_intrVec_8 = decoder2_io_out_bits_cf_intrVec_8; // @[src/main/scala/nutcore/frontend/IDU.scala 211:13]
  assign io_out_1_bits_cf_intrVec_9 = decoder2_io_out_bits_cf_intrVec_9; // @[src/main/scala/nutcore/frontend/IDU.scala 211:13]
  assign io_out_1_bits_cf_intrVec_10 = decoder2_io_out_bits_cf_intrVec_10; // @[src/main/scala/nutcore/frontend/IDU.scala 211:13]
  assign io_out_1_bits_cf_intrVec_11 = decoder2_io_out_bits_cf_intrVec_11; // @[src/main/scala/nutcore/frontend/IDU.scala 211:13]
  assign decoder1_io_in_valid = io_in_0_valid; // @[src/main/scala/nutcore/frontend/IDU.scala 208:12]
  assign decoder1_io_in_bits_instr = io_in_0_bits_instr; // @[src/main/scala/nutcore/frontend/IDU.scala 208:12]
  assign decoder1_io_in_bits_pc = io_in_0_bits_pc; // @[src/main/scala/nutcore/frontend/IDU.scala 208:12]
  assign decoder1_io_in_bits_pnpc = io_in_0_bits_pnpc; // @[src/main/scala/nutcore/frontend/IDU.scala 208:12]
  assign decoder1_io_in_bits_brIdx = io_in_0_bits_brIdx; // @[src/main/scala/nutcore/frontend/IDU.scala 208:12]
  assign decoder1_io_out_ready = io_out_0_ready; // @[src/main/scala/nutcore/frontend/IDU.scala 210:13]
  assign decoder1_intrVecIDU = intrVec;
  assign decoder2_intrVecIDU = intrVec;
endmodule
module FlushableQueue(
  input         clock,
  input         reset,
  output        io_enq_ready, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  input         io_enq_valid, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  input  [63:0] io_enq_bits_instr, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  input  [38:0] io_enq_bits_pc, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  input  [38:0] io_enq_bits_pnpc, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  input  [3:0]  io_enq_bits_brIdx, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  input         io_deq_ready, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_valid, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output [63:0] io_deq_bits_instr, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output [38:0] io_deq_bits_pc, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output [38:0] io_deq_bits_pnpc, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output [3:0]  io_deq_bits_brIdx, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  input         io_flush // @[src/main/scala/utils/FlushableQueue.scala 21:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] regs_0_instr; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [38:0] regs_0_pc; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [38:0] regs_0_pnpc; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [3:0] regs_0_brIdx; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [63:0] regs_1_instr; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [38:0] regs_1_pc; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [38:0] regs_1_pnpc; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [3:0] regs_1_brIdx; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [63:0] regs_2_instr; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [38:0] regs_2_pc; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [38:0] regs_2_pnpc; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [3:0] regs_2_brIdx; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [63:0] regs_3_instr; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [38:0] regs_3_pc; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [38:0] regs_3_pnpc; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [3:0] regs_3_brIdx; // @[src/main/scala/utils/RegMem.scala 7:21]
  reg [1:0] enq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg [1:0] deq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  maybe_full; // @[src/main/scala/utils/FlushableQueue.scala 26:35]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[src/main/scala/utils/FlushableQueue.scala 28:41]
  wire  empty = ptr_match & ~maybe_full; // @[src/main/scala/utils/FlushableQueue.scala 29:33]
  wire  full = ptr_match & maybe_full; // @[src/main/scala/utils/FlushableQueue.scala 30:32]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [1:0] _value_T_1 = enq_ptr_value + 2'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire [1:0] _value_T_3 = deq_ptr_value + 2'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire [63:0] _GEN_316 = 2'h1 == deq_ptr_value ? regs_1_instr : regs_0_instr; // @[src/main/scala/utils/FlushableQueue.scala 47:{15,15}]
  wire [63:0] _GEN_317 = 2'h2 == deq_ptr_value ? regs_2_instr : _GEN_316; // @[src/main/scala/utils/FlushableQueue.scala 47:{15,15}]
  wire [38:0] _GEN_320 = 2'h1 == deq_ptr_value ? regs_1_pc : regs_0_pc; // @[src/main/scala/utils/FlushableQueue.scala 47:{15,15}]
  wire [38:0] _GEN_321 = 2'h2 == deq_ptr_value ? regs_2_pc : _GEN_320; // @[src/main/scala/utils/FlushableQueue.scala 47:{15,15}]
  wire [38:0] _GEN_324 = 2'h1 == deq_ptr_value ? regs_1_pnpc : regs_0_pnpc; // @[src/main/scala/utils/FlushableQueue.scala 47:{15,15}]
  wire [38:0] _GEN_325 = 2'h2 == deq_ptr_value ? regs_2_pnpc : _GEN_324; // @[src/main/scala/utils/FlushableQueue.scala 47:{15,15}]
  wire [3:0] _GEN_452 = 2'h1 == deq_ptr_value ? regs_1_brIdx : regs_0_brIdx; // @[src/main/scala/utils/FlushableQueue.scala 47:{15,15}]
  wire [3:0] _GEN_453 = 2'h2 == deq_ptr_value ? regs_2_brIdx : _GEN_452; // @[src/main/scala/utils/FlushableQueue.scala 47:{15,15}]
  assign io_enq_ready = ~full; // @[src/main/scala/utils/FlushableQueue.scala 46:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/utils/FlushableQueue.scala 45:19]
  assign io_deq_bits_instr = 2'h3 == deq_ptr_value ? regs_3_instr : _GEN_317; // @[src/main/scala/utils/FlushableQueue.scala 47:{15,15}]
  assign io_deq_bits_pc = 2'h3 == deq_ptr_value ? regs_3_pc : _GEN_321; // @[src/main/scala/utils/FlushableQueue.scala 47:{15,15}]
  assign io_deq_bits_pnpc = 2'h3 == deq_ptr_value ? regs_3_pnpc : _GEN_325; // @[src/main/scala/utils/FlushableQueue.scala 47:{15,15}]
  assign io_deq_bits_brIdx = 2'h3 == deq_ptr_value ? regs_3_brIdx : _GEN_453; // @[src/main/scala/utils/FlushableQueue.scala 47:{15,15}]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_0_instr <= 64'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (do_enq) begin // @[src/main/scala/utils/FlushableQueue.scala 34:17]
      if (2'h0 == enq_ptr_value) begin // @[src/main/scala/utils/FlushableQueue.scala 35:24]
        regs_0_instr <= io_enq_bits_instr; // @[src/main/scala/utils/FlushableQueue.scala 35:24]
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_0_pc <= 39'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (do_enq) begin // @[src/main/scala/utils/FlushableQueue.scala 34:17]
      if (2'h0 == enq_ptr_value) begin // @[src/main/scala/utils/FlushableQueue.scala 35:24]
        regs_0_pc <= io_enq_bits_pc; // @[src/main/scala/utils/FlushableQueue.scala 35:24]
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_0_pnpc <= 39'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (do_enq) begin // @[src/main/scala/utils/FlushableQueue.scala 34:17]
      if (2'h0 == enq_ptr_value) begin // @[src/main/scala/utils/FlushableQueue.scala 35:24]
        regs_0_pnpc <= io_enq_bits_pnpc; // @[src/main/scala/utils/FlushableQueue.scala 35:24]
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_0_brIdx <= 4'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (do_enq) begin // @[src/main/scala/utils/FlushableQueue.scala 34:17]
      if (2'h0 == enq_ptr_value) begin // @[src/main/scala/utils/FlushableQueue.scala 35:24]
        regs_0_brIdx <= io_enq_bits_brIdx; // @[src/main/scala/utils/FlushableQueue.scala 35:24]
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_1_instr <= 64'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (do_enq) begin // @[src/main/scala/utils/FlushableQueue.scala 34:17]
      if (2'h1 == enq_ptr_value) begin // @[src/main/scala/utils/FlushableQueue.scala 35:24]
        regs_1_instr <= io_enq_bits_instr; // @[src/main/scala/utils/FlushableQueue.scala 35:24]
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_1_pc <= 39'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (do_enq) begin // @[src/main/scala/utils/FlushableQueue.scala 34:17]
      if (2'h1 == enq_ptr_value) begin // @[src/main/scala/utils/FlushableQueue.scala 35:24]
        regs_1_pc <= io_enq_bits_pc; // @[src/main/scala/utils/FlushableQueue.scala 35:24]
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_1_pnpc <= 39'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (do_enq) begin // @[src/main/scala/utils/FlushableQueue.scala 34:17]
      if (2'h1 == enq_ptr_value) begin // @[src/main/scala/utils/FlushableQueue.scala 35:24]
        regs_1_pnpc <= io_enq_bits_pnpc; // @[src/main/scala/utils/FlushableQueue.scala 35:24]
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_1_brIdx <= 4'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (do_enq) begin // @[src/main/scala/utils/FlushableQueue.scala 34:17]
      if (2'h1 == enq_ptr_value) begin // @[src/main/scala/utils/FlushableQueue.scala 35:24]
        regs_1_brIdx <= io_enq_bits_brIdx; // @[src/main/scala/utils/FlushableQueue.scala 35:24]
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_2_instr <= 64'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (do_enq) begin // @[src/main/scala/utils/FlushableQueue.scala 34:17]
      if (2'h2 == enq_ptr_value) begin // @[src/main/scala/utils/FlushableQueue.scala 35:24]
        regs_2_instr <= io_enq_bits_instr; // @[src/main/scala/utils/FlushableQueue.scala 35:24]
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_2_pc <= 39'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (do_enq) begin // @[src/main/scala/utils/FlushableQueue.scala 34:17]
      if (2'h2 == enq_ptr_value) begin // @[src/main/scala/utils/FlushableQueue.scala 35:24]
        regs_2_pc <= io_enq_bits_pc; // @[src/main/scala/utils/FlushableQueue.scala 35:24]
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_2_pnpc <= 39'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (do_enq) begin // @[src/main/scala/utils/FlushableQueue.scala 34:17]
      if (2'h2 == enq_ptr_value) begin // @[src/main/scala/utils/FlushableQueue.scala 35:24]
        regs_2_pnpc <= io_enq_bits_pnpc; // @[src/main/scala/utils/FlushableQueue.scala 35:24]
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_2_brIdx <= 4'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (do_enq) begin // @[src/main/scala/utils/FlushableQueue.scala 34:17]
      if (2'h2 == enq_ptr_value) begin // @[src/main/scala/utils/FlushableQueue.scala 35:24]
        regs_2_brIdx <= io_enq_bits_brIdx; // @[src/main/scala/utils/FlushableQueue.scala 35:24]
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_3_instr <= 64'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (do_enq) begin // @[src/main/scala/utils/FlushableQueue.scala 34:17]
      if (2'h3 == enq_ptr_value) begin // @[src/main/scala/utils/FlushableQueue.scala 35:24]
        regs_3_instr <= io_enq_bits_instr; // @[src/main/scala/utils/FlushableQueue.scala 35:24]
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_3_pc <= 39'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (do_enq) begin // @[src/main/scala/utils/FlushableQueue.scala 34:17]
      if (2'h3 == enq_ptr_value) begin // @[src/main/scala/utils/FlushableQueue.scala 35:24]
        regs_3_pc <= io_enq_bits_pc; // @[src/main/scala/utils/FlushableQueue.scala 35:24]
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_3_pnpc <= 39'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (do_enq) begin // @[src/main/scala/utils/FlushableQueue.scala 34:17]
      if (2'h3 == enq_ptr_value) begin // @[src/main/scala/utils/FlushableQueue.scala 35:24]
        regs_3_pnpc <= io_enq_bits_pnpc; // @[src/main/scala/utils/FlushableQueue.scala 35:24]
      end
    end
    if (reset) begin // @[src/main/scala/utils/RegMem.scala 7:21]
      regs_3_brIdx <= 4'h0; // @[src/main/scala/utils/RegMem.scala 7:21]
    end else if (do_enq) begin // @[src/main/scala/utils/FlushableQueue.scala 34:17]
      if (2'h3 == enq_ptr_value) begin // @[src/main/scala/utils/FlushableQueue.scala 35:24]
        regs_3_brIdx <= io_enq_bits_brIdx; // @[src/main/scala/utils/FlushableQueue.scala 35:24]
      end
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      enq_ptr_value <= 2'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (io_flush) begin // @[src/main/scala/utils/FlushableQueue.scala 62:19]
      enq_ptr_value <= 2'h0; // @[src/main/scala/utils/FlushableQueue.scala 64:21]
    end else if (do_enq) begin // @[src/main/scala/utils/FlushableQueue.scala 34:17]
      enq_ptr_value <= _value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      deq_ptr_value <= 2'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (io_flush) begin // @[src/main/scala/utils/FlushableQueue.scala 62:19]
      deq_ptr_value <= 2'h0; // @[src/main/scala/utils/FlushableQueue.scala 65:21]
    end else if (do_deq) begin // @[src/main/scala/utils/FlushableQueue.scala 38:17]
      deq_ptr_value <= _value_T_3; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/utils/FlushableQueue.scala 26:35]
      maybe_full <= 1'h0; // @[src/main/scala/utils/FlushableQueue.scala 26:35]
    end else if (io_flush) begin // @[src/main/scala/utils/FlushableQueue.scala 62:19]
      maybe_full <= 1'h0; // @[src/main/scala/utils/FlushableQueue.scala 67:16]
    end else if (do_enq != do_deq) begin // @[src/main/scala/utils/FlushableQueue.scala 41:28]
      maybe_full <= do_enq; // @[src/main/scala/utils/FlushableQueue.scala 42:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  regs_0_instr = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  regs_0_pc = _RAND_1[38:0];
  _RAND_2 = {2{`RANDOM}};
  regs_0_pnpc = _RAND_2[38:0];
  _RAND_3 = {1{`RANDOM}};
  regs_0_brIdx = _RAND_3[3:0];
  _RAND_4 = {2{`RANDOM}};
  regs_1_instr = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  regs_1_pc = _RAND_5[38:0];
  _RAND_6 = {2{`RANDOM}};
  regs_1_pnpc = _RAND_6[38:0];
  _RAND_7 = {1{`RANDOM}};
  regs_1_brIdx = _RAND_7[3:0];
  _RAND_8 = {2{`RANDOM}};
  regs_2_instr = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  regs_2_pc = _RAND_9[38:0];
  _RAND_10 = {2{`RANDOM}};
  regs_2_pnpc = _RAND_10[38:0];
  _RAND_11 = {1{`RANDOM}};
  regs_2_brIdx = _RAND_11[3:0];
  _RAND_12 = {2{`RANDOM}};
  regs_3_instr = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  regs_3_pc = _RAND_13[38:0];
  _RAND_14 = {2{`RANDOM}};
  regs_3_pnpc = _RAND_14[38:0];
  _RAND_15 = {1{`RANDOM}};
  regs_3_brIdx = _RAND_15[3:0];
  _RAND_16 = {1{`RANDOM}};
  enq_ptr_value = _RAND_16[1:0];
  _RAND_17 = {1{`RANDOM}};
  deq_ptr_value = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  maybe_full = _RAND_18[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Frontend_inorder(
  input         clock,
  input         reset,
  input         io_imem_req_ready, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output        io_imem_req_valid, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output [38:0] io_imem_req_bits_addr, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output [86:0] io_imem_req_bits_user, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output        io_imem_resp_ready, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  input         io_imem_resp_valid, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  input  [63:0] io_imem_resp_bits_rdata, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  input  [86:0] io_imem_resp_bits_user, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  input         io_out_0_ready, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output        io_out_0_valid, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output [63:0] io_out_0_bits_cf_instr, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output [38:0] io_out_0_bits_cf_pc, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output [38:0] io_out_0_bits_cf_pnpc, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output        io_out_0_bits_cf_exceptionVec_1, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output        io_out_0_bits_cf_exceptionVec_2, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output        io_out_0_bits_cf_intrVec_0, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output        io_out_0_bits_cf_intrVec_1, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output        io_out_0_bits_cf_intrVec_2, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output        io_out_0_bits_cf_intrVec_3, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output        io_out_0_bits_cf_intrVec_4, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output        io_out_0_bits_cf_intrVec_5, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output        io_out_0_bits_cf_intrVec_6, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output        io_out_0_bits_cf_intrVec_7, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output        io_out_0_bits_cf_intrVec_8, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output        io_out_0_bits_cf_intrVec_9, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output        io_out_0_bits_cf_intrVec_10, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output        io_out_0_bits_cf_intrVec_11, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output [3:0]  io_out_0_bits_cf_brIdx, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output        io_out_0_bits_ctrl_src1Type, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output        io_out_0_bits_ctrl_src2Type, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output [2:0]  io_out_0_bits_ctrl_fuType, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output [6:0]  io_out_0_bits_ctrl_fuOpType, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output [4:0]  io_out_0_bits_ctrl_rfSrc1, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output [4:0]  io_out_0_bits_ctrl_rfSrc2, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output        io_out_0_bits_ctrl_rfWen, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output [4:0]  io_out_0_bits_ctrl_rfDest, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output [63:0] io_out_0_bits_data_imm, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output        io_out_1_bits_cf_intrVec_0, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output        io_out_1_bits_cf_intrVec_1, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output        io_out_1_bits_cf_intrVec_2, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output        io_out_1_bits_cf_intrVec_3, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output        io_out_1_bits_cf_intrVec_4, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output        io_out_1_bits_cf_intrVec_5, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output        io_out_1_bits_cf_intrVec_6, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output        io_out_1_bits_cf_intrVec_7, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output        io_out_1_bits_cf_intrVec_8, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output        io_out_1_bits_cf_intrVec_9, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output        io_out_1_bits_cf_intrVec_10, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output        io_out_1_bits_cf_intrVec_11, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  output [3:0]  io_flushVec, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  input  [38:0] io_redirect_target, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  input         io_redirect_valid, // @[src/main/scala/nutcore/frontend/Frontend.scala 40:14]
  input         flushICache,
  input         REG_valid,
  input  [38:0] REG_pc,
  input         REG_isMissPredict,
  input  [38:0] REG_actualTarget,
  input         REG_actualTaken,
  input  [6:0]  REG_fuOpType,
  input  [1:0]  REG_btbType,
  input         REG_isRVC,
  input  [11:0] intrVec,
  input         flushTLB
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  ifu_clock; // @[src/main/scala/nutcore/frontend/Frontend.scala 98:20]
  wire  ifu_reset; // @[src/main/scala/nutcore/frontend/Frontend.scala 98:20]
  wire  ifu_io_imem_req_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 98:20]
  wire  ifu_io_imem_req_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 98:20]
  wire [38:0] ifu_io_imem_req_bits_addr; // @[src/main/scala/nutcore/frontend/Frontend.scala 98:20]
  wire [81:0] ifu_io_imem_req_bits_user; // @[src/main/scala/nutcore/frontend/Frontend.scala 98:20]
  wire  ifu_io_imem_resp_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 98:20]
  wire  ifu_io_imem_resp_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 98:20]
  wire [63:0] ifu_io_imem_resp_bits_rdata; // @[src/main/scala/nutcore/frontend/Frontend.scala 98:20]
  wire [81:0] ifu_io_imem_resp_bits_user; // @[src/main/scala/nutcore/frontend/Frontend.scala 98:20]
  wire  ifu_io_out_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 98:20]
  wire  ifu_io_out_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 98:20]
  wire [63:0] ifu_io_out_bits_instr; // @[src/main/scala/nutcore/frontend/Frontend.scala 98:20]
  wire [38:0] ifu_io_out_bits_pc; // @[src/main/scala/nutcore/frontend/Frontend.scala 98:20]
  wire [38:0] ifu_io_out_bits_pnpc; // @[src/main/scala/nutcore/frontend/Frontend.scala 98:20]
  wire [3:0] ifu_io_out_bits_brIdx; // @[src/main/scala/nutcore/frontend/Frontend.scala 98:20]
  wire [38:0] ifu_io_redirect_target; // @[src/main/scala/nutcore/frontend/Frontend.scala 98:20]
  wire  ifu_io_redirect_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 98:20]
  wire [3:0] ifu_io_flushVec; // @[src/main/scala/nutcore/frontend/Frontend.scala 98:20]
  wire  ifu_flushICache; // @[src/main/scala/nutcore/frontend/Frontend.scala 98:20]
  wire  ifu_REG_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 98:20]
  wire [38:0] ifu_REG_pc; // @[src/main/scala/nutcore/frontend/Frontend.scala 98:20]
  wire  ifu_REG_isMissPredict; // @[src/main/scala/nutcore/frontend/Frontend.scala 98:20]
  wire [38:0] ifu_REG_actualTarget; // @[src/main/scala/nutcore/frontend/Frontend.scala 98:20]
  wire  ifu_REG_actualTaken; // @[src/main/scala/nutcore/frontend/Frontend.scala 98:20]
  wire [6:0] ifu_REG_fuOpType; // @[src/main/scala/nutcore/frontend/Frontend.scala 98:20]
  wire [1:0] ifu_REG_btbType; // @[src/main/scala/nutcore/frontend/Frontend.scala 98:20]
  wire  ifu_REG_isRVC; // @[src/main/scala/nutcore/frontend/Frontend.scala 98:20]
  wire  ifu_flushTLB; // @[src/main/scala/nutcore/frontend/Frontend.scala 98:20]
  wire  ibf_clock; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:19]
  wire  ibf_reset; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:19]
  wire  ibf_io_in_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:19]
  wire  ibf_io_in_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:19]
  wire [63:0] ibf_io_in_bits_instr; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:19]
  wire [38:0] ibf_io_in_bits_pc; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:19]
  wire [38:0] ibf_io_in_bits_pnpc; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:19]
  wire [3:0] ibf_io_in_bits_brIdx; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:19]
  wire  ibf_io_out_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:19]
  wire  ibf_io_out_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:19]
  wire [63:0] ibf_io_out_bits_instr; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:19]
  wire [38:0] ibf_io_out_bits_pc; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:19]
  wire [38:0] ibf_io_out_bits_pnpc; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:19]
  wire [3:0] ibf_io_out_bits_brIdx; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:19]
  wire  ibf_io_flush; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:19]
  wire  idu_io_in_0_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire  idu_io_in_0_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire [63:0] idu_io_in_0_bits_instr; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire [38:0] idu_io_in_0_bits_pc; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire [38:0] idu_io_in_0_bits_pnpc; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire [3:0] idu_io_in_0_bits_brIdx; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire  idu_io_out_0_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire  idu_io_out_0_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire [63:0] idu_io_out_0_bits_cf_instr; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire [38:0] idu_io_out_0_bits_cf_pc; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire [38:0] idu_io_out_0_bits_cf_pnpc; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire  idu_io_out_0_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire  idu_io_out_0_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire  idu_io_out_0_bits_cf_intrVec_0; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire  idu_io_out_0_bits_cf_intrVec_1; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire  idu_io_out_0_bits_cf_intrVec_2; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire  idu_io_out_0_bits_cf_intrVec_3; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire  idu_io_out_0_bits_cf_intrVec_4; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire  idu_io_out_0_bits_cf_intrVec_5; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire  idu_io_out_0_bits_cf_intrVec_6; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire  idu_io_out_0_bits_cf_intrVec_7; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire  idu_io_out_0_bits_cf_intrVec_8; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire  idu_io_out_0_bits_cf_intrVec_9; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire  idu_io_out_0_bits_cf_intrVec_10; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire  idu_io_out_0_bits_cf_intrVec_11; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire [3:0] idu_io_out_0_bits_cf_brIdx; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire  idu_io_out_0_bits_ctrl_src1Type; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire  idu_io_out_0_bits_ctrl_src2Type; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire [2:0] idu_io_out_0_bits_ctrl_fuType; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire [6:0] idu_io_out_0_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire [4:0] idu_io_out_0_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire [4:0] idu_io_out_0_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire  idu_io_out_0_bits_ctrl_rfWen; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire [4:0] idu_io_out_0_bits_ctrl_rfDest; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire [63:0] idu_io_out_0_bits_data_imm; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire  idu_io_out_1_bits_cf_intrVec_0; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire  idu_io_out_1_bits_cf_intrVec_1; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire  idu_io_out_1_bits_cf_intrVec_2; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire  idu_io_out_1_bits_cf_intrVec_3; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire  idu_io_out_1_bits_cf_intrVec_4; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire  idu_io_out_1_bits_cf_intrVec_5; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire  idu_io_out_1_bits_cf_intrVec_6; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire  idu_io_out_1_bits_cf_intrVec_7; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire  idu_io_out_1_bits_cf_intrVec_8; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire  idu_io_out_1_bits_cf_intrVec_9; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire  idu_io_out_1_bits_cf_intrVec_10; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire  idu_io_out_1_bits_cf_intrVec_11; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire [11:0] idu_intrVec; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
  wire  ibf_io_in_q_clock; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_reset; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_enq_ready; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_enq_valid; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire [63:0] ibf_io_in_q_io_enq_bits_instr; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire [38:0] ibf_io_in_q_io_enq_bits_pc; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire [38:0] ibf_io_in_q_io_enq_bits_pnpc; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire [3:0] ibf_io_in_q_io_enq_bits_brIdx; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_ready; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_valid; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire [63:0] ibf_io_in_q_io_deq_bits_instr; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire [38:0] ibf_io_in_q_io_deq_bits_pc; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire [38:0] ibf_io_in_q_io_deq_bits_pnpc; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire [3:0] ibf_io_in_q_io_deq_bits_brIdx; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_flush; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  _T_1 = idu_io_out_0_ready & idu_io_out_0_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  valid; // @[src/main/scala/utils/Pipeline.scala 24:24]
  wire  _GEN_0 = _T_1 ? 1'h0 : valid; // @[src/main/scala/utils/Pipeline.scala 24:24 25:{25,33}]
  wire  _T_3 = ibf_io_out_valid & idu_io_in_0_ready; // @[src/main/scala/utils/Pipeline.scala 26:22]
  wire  _GEN_1 = ibf_io_out_valid & idu_io_in_0_ready | _GEN_0; // @[src/main/scala/utils/Pipeline.scala 26:{38,46}]
  reg [63:0] idu_io_in_0_bits_r_instr; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [38:0] idu_io_in_0_bits_r_pc; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [38:0] idu_io_in_0_bits_r_pnpc; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [3:0] idu_io_in_0_bits_r_brIdx; // @[src/main/scala/utils/Pipeline.scala 30:28]
  IFU_inorder ifu ( // @[src/main/scala/nutcore/frontend/Frontend.scala 98:20]
    .clock(ifu_clock),
    .reset(ifu_reset),
    .io_imem_req_ready(ifu_io_imem_req_ready),
    .io_imem_req_valid(ifu_io_imem_req_valid),
    .io_imem_req_bits_addr(ifu_io_imem_req_bits_addr),
    .io_imem_req_bits_user(ifu_io_imem_req_bits_user),
    .io_imem_resp_ready(ifu_io_imem_resp_ready),
    .io_imem_resp_valid(ifu_io_imem_resp_valid),
    .io_imem_resp_bits_rdata(ifu_io_imem_resp_bits_rdata),
    .io_imem_resp_bits_user(ifu_io_imem_resp_bits_user),
    .io_out_ready(ifu_io_out_ready),
    .io_out_valid(ifu_io_out_valid),
    .io_out_bits_instr(ifu_io_out_bits_instr),
    .io_out_bits_pc(ifu_io_out_bits_pc),
    .io_out_bits_pnpc(ifu_io_out_bits_pnpc),
    .io_out_bits_brIdx(ifu_io_out_bits_brIdx),
    .io_redirect_target(ifu_io_redirect_target),
    .io_redirect_valid(ifu_io_redirect_valid),
    .io_flushVec(ifu_io_flushVec),
    .flushICache(ifu_flushICache),
    .REG_valid(ifu_REG_valid),
    .REG_pc(ifu_REG_pc),
    .REG_isMissPredict(ifu_REG_isMissPredict),
    .REG_actualTarget(ifu_REG_actualTarget),
    .REG_actualTaken(ifu_REG_actualTaken),
    .REG_fuOpType(ifu_REG_fuOpType),
    .REG_btbType(ifu_REG_btbType),
    .REG_isRVC(ifu_REG_isRVC),
    .flushTLB(ifu_flushTLB)
  );
  NaiveRVCAlignBuffer ibf ( // @[src/main/scala/nutcore/frontend/Frontend.scala 99:19]
    .clock(ibf_clock),
    .reset(ibf_reset),
    .io_in_ready(ibf_io_in_ready),
    .io_in_valid(ibf_io_in_valid),
    .io_in_bits_instr(ibf_io_in_bits_instr),
    .io_in_bits_pc(ibf_io_in_bits_pc),
    .io_in_bits_pnpc(ibf_io_in_bits_pnpc),
    .io_in_bits_brIdx(ibf_io_in_bits_brIdx),
    .io_out_ready(ibf_io_out_ready),
    .io_out_valid(ibf_io_out_valid),
    .io_out_bits_instr(ibf_io_out_bits_instr),
    .io_out_bits_pc(ibf_io_out_bits_pc),
    .io_out_bits_pnpc(ibf_io_out_bits_pnpc),
    .io_out_bits_brIdx(ibf_io_out_bits_brIdx),
    .io_flush(ibf_io_flush)
  );
  IDU idu ( // @[src/main/scala/nutcore/frontend/Frontend.scala 100:20]
    .io_in_0_ready(idu_io_in_0_ready),
    .io_in_0_valid(idu_io_in_0_valid),
    .io_in_0_bits_instr(idu_io_in_0_bits_instr),
    .io_in_0_bits_pc(idu_io_in_0_bits_pc),
    .io_in_0_bits_pnpc(idu_io_in_0_bits_pnpc),
    .io_in_0_bits_brIdx(idu_io_in_0_bits_brIdx),
    .io_out_0_ready(idu_io_out_0_ready),
    .io_out_0_valid(idu_io_out_0_valid),
    .io_out_0_bits_cf_instr(idu_io_out_0_bits_cf_instr),
    .io_out_0_bits_cf_pc(idu_io_out_0_bits_cf_pc),
    .io_out_0_bits_cf_pnpc(idu_io_out_0_bits_cf_pnpc),
    .io_out_0_bits_cf_exceptionVec_1(idu_io_out_0_bits_cf_exceptionVec_1),
    .io_out_0_bits_cf_exceptionVec_2(idu_io_out_0_bits_cf_exceptionVec_2),
    .io_out_0_bits_cf_intrVec_0(idu_io_out_0_bits_cf_intrVec_0),
    .io_out_0_bits_cf_intrVec_1(idu_io_out_0_bits_cf_intrVec_1),
    .io_out_0_bits_cf_intrVec_2(idu_io_out_0_bits_cf_intrVec_2),
    .io_out_0_bits_cf_intrVec_3(idu_io_out_0_bits_cf_intrVec_3),
    .io_out_0_bits_cf_intrVec_4(idu_io_out_0_bits_cf_intrVec_4),
    .io_out_0_bits_cf_intrVec_5(idu_io_out_0_bits_cf_intrVec_5),
    .io_out_0_bits_cf_intrVec_6(idu_io_out_0_bits_cf_intrVec_6),
    .io_out_0_bits_cf_intrVec_7(idu_io_out_0_bits_cf_intrVec_7),
    .io_out_0_bits_cf_intrVec_8(idu_io_out_0_bits_cf_intrVec_8),
    .io_out_0_bits_cf_intrVec_9(idu_io_out_0_bits_cf_intrVec_9),
    .io_out_0_bits_cf_intrVec_10(idu_io_out_0_bits_cf_intrVec_10),
    .io_out_0_bits_cf_intrVec_11(idu_io_out_0_bits_cf_intrVec_11),
    .io_out_0_bits_cf_brIdx(idu_io_out_0_bits_cf_brIdx),
    .io_out_0_bits_ctrl_src1Type(idu_io_out_0_bits_ctrl_src1Type),
    .io_out_0_bits_ctrl_src2Type(idu_io_out_0_bits_ctrl_src2Type),
    .io_out_0_bits_ctrl_fuType(idu_io_out_0_bits_ctrl_fuType),
    .io_out_0_bits_ctrl_fuOpType(idu_io_out_0_bits_ctrl_fuOpType),
    .io_out_0_bits_ctrl_rfSrc1(idu_io_out_0_bits_ctrl_rfSrc1),
    .io_out_0_bits_ctrl_rfSrc2(idu_io_out_0_bits_ctrl_rfSrc2),
    .io_out_0_bits_ctrl_rfWen(idu_io_out_0_bits_ctrl_rfWen),
    .io_out_0_bits_ctrl_rfDest(idu_io_out_0_bits_ctrl_rfDest),
    .io_out_0_bits_data_imm(idu_io_out_0_bits_data_imm),
    .io_out_1_bits_cf_intrVec_0(idu_io_out_1_bits_cf_intrVec_0),
    .io_out_1_bits_cf_intrVec_1(idu_io_out_1_bits_cf_intrVec_1),
    .io_out_1_bits_cf_intrVec_2(idu_io_out_1_bits_cf_intrVec_2),
    .io_out_1_bits_cf_intrVec_3(idu_io_out_1_bits_cf_intrVec_3),
    .io_out_1_bits_cf_intrVec_4(idu_io_out_1_bits_cf_intrVec_4),
    .io_out_1_bits_cf_intrVec_5(idu_io_out_1_bits_cf_intrVec_5),
    .io_out_1_bits_cf_intrVec_6(idu_io_out_1_bits_cf_intrVec_6),
    .io_out_1_bits_cf_intrVec_7(idu_io_out_1_bits_cf_intrVec_7),
    .io_out_1_bits_cf_intrVec_8(idu_io_out_1_bits_cf_intrVec_8),
    .io_out_1_bits_cf_intrVec_9(idu_io_out_1_bits_cf_intrVec_9),
    .io_out_1_bits_cf_intrVec_10(idu_io_out_1_bits_cf_intrVec_10),
    .io_out_1_bits_cf_intrVec_11(idu_io_out_1_bits_cf_intrVec_11),
    .intrVec(idu_intrVec)
  );
  FlushableQueue ibf_io_in_q ( // @[src/main/scala/utils/FlushableQueue.scala 94:21]
    .clock(ibf_io_in_q_clock),
    .reset(ibf_io_in_q_reset),
    .io_enq_ready(ibf_io_in_q_io_enq_ready),
    .io_enq_valid(ibf_io_in_q_io_enq_valid),
    .io_enq_bits_instr(ibf_io_in_q_io_enq_bits_instr),
    .io_enq_bits_pc(ibf_io_in_q_io_enq_bits_pc),
    .io_enq_bits_pnpc(ibf_io_in_q_io_enq_bits_pnpc),
    .io_enq_bits_brIdx(ibf_io_in_q_io_enq_bits_brIdx),
    .io_deq_ready(ibf_io_in_q_io_deq_ready),
    .io_deq_valid(ibf_io_in_q_io_deq_valid),
    .io_deq_bits_instr(ibf_io_in_q_io_deq_bits_instr),
    .io_deq_bits_pc(ibf_io_in_q_io_deq_bits_pc),
    .io_deq_bits_pnpc(ibf_io_in_q_io_deq_bits_pnpc),
    .io_deq_bits_brIdx(ibf_io_in_q_io_deq_bits_brIdx),
    .io_flush(ibf_io_in_q_io_flush)
  );
  assign io_imem_req_valid = ifu_io_imem_req_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 119:11]
  assign io_imem_req_bits_addr = ifu_io_imem_req_bits_addr; // @[src/main/scala/nutcore/frontend/Frontend.scala 119:11]
  assign io_imem_req_bits_user = {{5'd0}, ifu_io_imem_req_bits_user}; // @[src/main/scala/nutcore/frontend/Frontend.scala 119:11]
  assign io_imem_resp_ready = ifu_io_imem_resp_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 119:11]
  assign io_out_0_valid = idu_io_out_0_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:10]
  assign io_out_0_bits_cf_instr = idu_io_out_0_bits_cf_instr; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:10]
  assign io_out_0_bits_cf_pc = idu_io_out_0_bits_cf_pc; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:10]
  assign io_out_0_bits_cf_pnpc = idu_io_out_0_bits_cf_pnpc; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:10]
  assign io_out_0_bits_cf_exceptionVec_1 = idu_io_out_0_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:10]
  assign io_out_0_bits_cf_exceptionVec_2 = idu_io_out_0_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:10]
  assign io_out_0_bits_cf_intrVec_0 = idu_io_out_0_bits_cf_intrVec_0; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:10]
  assign io_out_0_bits_cf_intrVec_1 = idu_io_out_0_bits_cf_intrVec_1; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:10]
  assign io_out_0_bits_cf_intrVec_2 = idu_io_out_0_bits_cf_intrVec_2; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:10]
  assign io_out_0_bits_cf_intrVec_3 = idu_io_out_0_bits_cf_intrVec_3; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:10]
  assign io_out_0_bits_cf_intrVec_4 = idu_io_out_0_bits_cf_intrVec_4; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:10]
  assign io_out_0_bits_cf_intrVec_5 = idu_io_out_0_bits_cf_intrVec_5; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:10]
  assign io_out_0_bits_cf_intrVec_6 = idu_io_out_0_bits_cf_intrVec_6; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:10]
  assign io_out_0_bits_cf_intrVec_7 = idu_io_out_0_bits_cf_intrVec_7; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:10]
  assign io_out_0_bits_cf_intrVec_8 = idu_io_out_0_bits_cf_intrVec_8; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:10]
  assign io_out_0_bits_cf_intrVec_9 = idu_io_out_0_bits_cf_intrVec_9; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:10]
  assign io_out_0_bits_cf_intrVec_10 = idu_io_out_0_bits_cf_intrVec_10; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:10]
  assign io_out_0_bits_cf_intrVec_11 = idu_io_out_0_bits_cf_intrVec_11; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:10]
  assign io_out_0_bits_cf_brIdx = idu_io_out_0_bits_cf_brIdx; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:10]
  assign io_out_0_bits_ctrl_src1Type = idu_io_out_0_bits_ctrl_src1Type; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:10]
  assign io_out_0_bits_ctrl_src2Type = idu_io_out_0_bits_ctrl_src2Type; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:10]
  assign io_out_0_bits_ctrl_fuType = idu_io_out_0_bits_ctrl_fuType; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:10]
  assign io_out_0_bits_ctrl_fuOpType = idu_io_out_0_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:10]
  assign io_out_0_bits_ctrl_rfSrc1 = idu_io_out_0_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:10]
  assign io_out_0_bits_ctrl_rfSrc2 = idu_io_out_0_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:10]
  assign io_out_0_bits_ctrl_rfWen = idu_io_out_0_bits_ctrl_rfWen; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:10]
  assign io_out_0_bits_ctrl_rfDest = idu_io_out_0_bits_ctrl_rfDest; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:10]
  assign io_out_0_bits_data_imm = idu_io_out_0_bits_data_imm; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:10]
  assign io_out_1_bits_cf_intrVec_0 = idu_io_out_1_bits_cf_intrVec_0; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:10]
  assign io_out_1_bits_cf_intrVec_1 = idu_io_out_1_bits_cf_intrVec_1; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:10]
  assign io_out_1_bits_cf_intrVec_2 = idu_io_out_1_bits_cf_intrVec_2; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:10]
  assign io_out_1_bits_cf_intrVec_3 = idu_io_out_1_bits_cf_intrVec_3; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:10]
  assign io_out_1_bits_cf_intrVec_4 = idu_io_out_1_bits_cf_intrVec_4; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:10]
  assign io_out_1_bits_cf_intrVec_5 = idu_io_out_1_bits_cf_intrVec_5; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:10]
  assign io_out_1_bits_cf_intrVec_6 = idu_io_out_1_bits_cf_intrVec_6; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:10]
  assign io_out_1_bits_cf_intrVec_7 = idu_io_out_1_bits_cf_intrVec_7; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:10]
  assign io_out_1_bits_cf_intrVec_8 = idu_io_out_1_bits_cf_intrVec_8; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:10]
  assign io_out_1_bits_cf_intrVec_9 = idu_io_out_1_bits_cf_intrVec_9; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:10]
  assign io_out_1_bits_cf_intrVec_10 = idu_io_out_1_bits_cf_intrVec_10; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:10]
  assign io_out_1_bits_cf_intrVec_11 = idu_io_out_1_bits_cf_intrVec_11; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:10]
  assign io_flushVec = ifu_io_flushVec; // @[src/main/scala/nutcore/frontend/Frontend.scala 116:15]
  assign ifu_clock = clock;
  assign ifu_reset = reset;
  assign ifu_io_imem_req_ready = io_imem_req_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 119:11]
  assign ifu_io_imem_resp_valid = io_imem_resp_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 119:11]
  assign ifu_io_imem_resp_bits_rdata = io_imem_resp_bits_rdata; // @[src/main/scala/nutcore/frontend/Frontend.scala 119:11]
  assign ifu_io_imem_resp_bits_user = io_imem_resp_bits_user[81:0]; // @[src/main/scala/nutcore/frontend/Frontend.scala 119:11]
  assign ifu_io_out_ready = ibf_io_in_q_io_enq_ready; // @[src/main/scala/utils/FlushableQueue.scala 98:17]
  assign ifu_io_redirect_target = io_redirect_target; // @[src/main/scala/nutcore/frontend/Frontend.scala 115:15]
  assign ifu_io_redirect_valid = io_redirect_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 115:15]
  assign ifu_flushICache = flushICache;
  assign ifu_REG_valid = REG_valid;
  assign ifu_REG_pc = REG_pc;
  assign ifu_REG_isMissPredict = REG_isMissPredict;
  assign ifu_REG_actualTarget = REG_actualTarget;
  assign ifu_REG_actualTaken = REG_actualTaken;
  assign ifu_REG_fuOpType = REG_fuOpType;
  assign ifu_REG_btbType = REG_btbType;
  assign ifu_REG_isRVC = REG_isRVC;
  assign ifu_flushTLB = flushTLB;
  assign ibf_clock = clock;
  assign ibf_reset = reset;
  assign ibf_io_in_valid = ibf_io_in_q_io_deq_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 106:11]
  assign ibf_io_in_bits_instr = ibf_io_in_q_io_deq_bits_instr; // @[src/main/scala/nutcore/frontend/Frontend.scala 106:11]
  assign ibf_io_in_bits_pc = ibf_io_in_q_io_deq_bits_pc; // @[src/main/scala/nutcore/frontend/Frontend.scala 106:11]
  assign ibf_io_in_bits_pnpc = ibf_io_in_q_io_deq_bits_pnpc; // @[src/main/scala/nutcore/frontend/Frontend.scala 106:11]
  assign ibf_io_in_bits_brIdx = ibf_io_in_q_io_deq_bits_brIdx; // @[src/main/scala/nutcore/frontend/Frontend.scala 106:11]
  assign ibf_io_out_ready = idu_io_in_0_ready; // @[src/main/scala/utils/Pipeline.scala 29:16]
  assign ibf_io_flush = ifu_io_flushVec[1]; // @[src/main/scala/nutcore/frontend/Frontend.scala 113:34]
  assign idu_io_in_0_valid = valid; // @[src/main/scala/utils/Pipeline.scala 31:17]
  assign idu_io_in_0_bits_instr = idu_io_in_0_bits_r_instr; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign idu_io_in_0_bits_pc = idu_io_in_0_bits_r_pc; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign idu_io_in_0_bits_pnpc = idu_io_in_0_bits_r_pnpc; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign idu_io_in_0_bits_brIdx = idu_io_in_0_bits_r_brIdx; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign idu_io_out_0_ready = io_out_0_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:10]
  assign idu_intrVec = intrVec;
  assign ibf_io_in_q_clock = clock;
  assign ibf_io_in_q_reset = reset;
  assign ibf_io_in_q_io_enq_valid = ifu_io_out_valid; // @[src/main/scala/utils/FlushableQueue.scala 95:22]
  assign ibf_io_in_q_io_enq_bits_instr = ifu_io_out_bits_instr; // @[src/main/scala/utils/FlushableQueue.scala 96:21]
  assign ibf_io_in_q_io_enq_bits_pc = ifu_io_out_bits_pc; // @[src/main/scala/utils/FlushableQueue.scala 96:21]
  assign ibf_io_in_q_io_enq_bits_pnpc = ifu_io_out_bits_pnpc; // @[src/main/scala/utils/FlushableQueue.scala 96:21]
  assign ibf_io_in_q_io_enq_bits_brIdx = ifu_io_out_bits_brIdx; // @[src/main/scala/utils/FlushableQueue.scala 96:21]
  assign ibf_io_in_q_io_deq_ready = ibf_io_in_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 106:11]
  assign ibf_io_in_q_io_flush = ifu_io_flushVec[0]; // @[src/main/scala/nutcore/frontend/Frontend.scala 109:58]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/Pipeline.scala 24:24]
      valid <= 1'h0; // @[src/main/scala/utils/Pipeline.scala 24:24]
    end else if (ifu_io_flushVec[1]) begin // @[src/main/scala/utils/Pipeline.scala 27:20]
      valid <= 1'h0; // @[src/main/scala/utils/Pipeline.scala 27:28]
    end else begin
      valid <= _GEN_1;
    end
    if (_T_3) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      idu_io_in_0_bits_r_instr <= ibf_io_out_bits_instr; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_3) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      idu_io_in_0_bits_r_pc <= ibf_io_out_bits_pc; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_3) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      idu_io_in_0_bits_r_pnpc <= ibf_io_out_bits_pnpc; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_3) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      idu_io_in_0_bits_r_brIdx <= ibf_io_out_bits_brIdx; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  valid = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  idu_io_in_0_bits_r_instr = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  idu_io_in_0_bits_r_pc = _RAND_2[38:0];
  _RAND_3 = {2{`RANDOM}};
  idu_io_in_0_bits_r_pnpc = _RAND_3[38:0];
  _RAND_4 = {1{`RANDOM}};
  idu_io_in_0_bits_r_brIdx = _RAND_4[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ISU(
  input         clock,
  input         reset,
  output        io_in_0_ready, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_valid, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [63:0] io_in_0_bits_cf_instr, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [38:0] io_in_0_bits_cf_pc, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [38:0] io_in_0_bits_cf_pnpc, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_exceptionVec_1, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_exceptionVec_2, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_intrVec_0, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_intrVec_1, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_intrVec_2, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_intrVec_3, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_intrVec_4, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_intrVec_5, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_intrVec_6, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_intrVec_7, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_intrVec_8, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_intrVec_9, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_intrVec_10, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_intrVec_11, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [3:0]  io_in_0_bits_cf_brIdx, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_ctrl_src1Type, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_ctrl_src2Type, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [2:0]  io_in_0_bits_ctrl_fuType, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [6:0]  io_in_0_bits_ctrl_fuOpType, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [4:0]  io_in_0_bits_ctrl_rfSrc1, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [4:0]  io_in_0_bits_ctrl_rfSrc2, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_ctrl_rfWen, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [4:0]  io_in_0_bits_ctrl_rfDest, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [63:0] io_in_0_bits_data_imm, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_out_ready, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_valid, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [63:0] io_out_bits_cf_instr, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [38:0] io_out_bits_cf_pc, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [38:0] io_out_bits_cf_pnpc, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_exceptionVec_1, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_exceptionVec_2, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_intrVec_0, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_intrVec_1, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_intrVec_2, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_intrVec_3, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_intrVec_4, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_intrVec_5, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_intrVec_6, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_intrVec_7, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_intrVec_8, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_intrVec_9, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_intrVec_10, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_intrVec_11, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [3:0]  io_out_bits_cf_brIdx, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [2:0]  io_out_bits_ctrl_fuType, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [6:0]  io_out_bits_ctrl_fuOpType, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [4:0]  io_out_bits_ctrl_rfSrc1, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [4:0]  io_out_bits_ctrl_rfSrc2, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_ctrl_rfWen, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [4:0]  io_out_bits_ctrl_rfDest, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [63:0] io_out_bits_data_src1, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [63:0] io_out_bits_data_src2, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [63:0] io_out_bits_data_imm, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_wb_rfWen, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [4:0]  io_wb_rfDest, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [63:0] io_wb_rfData, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_forward_valid, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_forward_wb_rfWen, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [4:0]  io_forward_wb_rfDest, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [63:0] io_forward_wb_rfData, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [2:0]  io_forward_fuType, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_flush // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
`endif // RANDOMIZE_REG_INIT
  wire  forwardRfWen = io_forward_wb_rfWen & io_forward_valid; // @[src/main/scala/nutcore/backend/seq/ISU.scala 43:42]
  wire  dontForward1 = io_forward_fuType != 3'h0 & io_forward_fuType != 3'h1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 44:57]
  wire  src1DependEX = io_in_0_bits_ctrl_rfSrc1 != 5'h0 & io_in_0_bits_ctrl_rfSrc1 == io_forward_wb_rfDest &
    forwardRfWen; // @[src/main/scala/nutcore/backend/seq/ISU.scala 41:100]
  wire  src2DependEX = io_in_0_bits_ctrl_rfSrc2 != 5'h0 & io_in_0_bits_ctrl_rfSrc2 == io_forward_wb_rfDest &
    forwardRfWen; // @[src/main/scala/nutcore/backend/seq/ISU.scala 41:100]
  wire  src1DependWB = io_in_0_bits_ctrl_rfSrc1 != 5'h0 & io_in_0_bits_ctrl_rfSrc1 == io_wb_rfDest & io_wb_rfWen; // @[src/main/scala/nutcore/backend/seq/ISU.scala 41:100]
  wire  src2DependWB = io_in_0_bits_ctrl_rfSrc2 != 5'h0 & io_in_0_bits_ctrl_rfSrc2 == io_wb_rfDest & io_wb_rfWen; // @[src/main/scala/nutcore/backend/seq/ISU.scala 41:100]
  wire  _src1ForwardNextCycle_T = ~dontForward1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 50:46]
  wire  src1ForwardNextCycle = src1DependEX & ~dontForward1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 50:43]
  wire  src2ForwardNextCycle = src2DependEX & _src1ForwardNextCycle_T; // @[src/main/scala/nutcore/backend/seq/ISU.scala 51:43]
  wire  _src1Forward_T_1 = dontForward1 ? ~src1DependEX : 1'h1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 52:40]
  wire  src1Forward = src1DependWB & _src1Forward_T_1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 52:34]
  wire  _src2Forward_T_1 = dontForward1 ? ~src2DependEX : 1'h1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 53:40]
  wire  src2Forward = src2DependWB & _src2Forward_T_1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 53:34]
  reg [31:0] busy; // @[src/main/scala/nutcore/RF.scala 50:21]
  wire [31:0] _src1Ready_T = busy >> io_in_0_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/RF.scala 51:37]
  wire  src1Ready = ~_src1Ready_T[0] | src1ForwardNextCycle | src1Forward; // @[src/main/scala/nutcore/backend/seq/ISU.scala 56:62]
  wire [31:0] _src2Ready_T = busy >> io_in_0_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/RF.scala 51:37]
  wire  src2Ready = ~_src2Ready_T[0] | src2ForwardNextCycle | src2Forward; // @[src/main/scala/nutcore/backend/seq/ISU.scala 57:62]
  reg [63:0] rf_0; // @[src/main/scala/nutcore/RF.scala 33:15]
  reg [63:0] rf_1; // @[src/main/scala/nutcore/RF.scala 33:15]
  reg [63:0] rf_2; // @[src/main/scala/nutcore/RF.scala 33:15]
  reg [63:0] rf_3; // @[src/main/scala/nutcore/RF.scala 33:15]
  reg [63:0] rf_4; // @[src/main/scala/nutcore/RF.scala 33:15]
  reg [63:0] rf_5; // @[src/main/scala/nutcore/RF.scala 33:15]
  reg [63:0] rf_6; // @[src/main/scala/nutcore/RF.scala 33:15]
  reg [63:0] rf_7; // @[src/main/scala/nutcore/RF.scala 33:15]
  reg [63:0] rf_8; // @[src/main/scala/nutcore/RF.scala 33:15]
  reg [63:0] rf_9; // @[src/main/scala/nutcore/RF.scala 33:15]
  reg [63:0] rf_10; // @[src/main/scala/nutcore/RF.scala 33:15]
  reg [63:0] rf_11; // @[src/main/scala/nutcore/RF.scala 33:15]
  reg [63:0] rf_12; // @[src/main/scala/nutcore/RF.scala 33:15]
  reg [63:0] rf_13; // @[src/main/scala/nutcore/RF.scala 33:15]
  reg [63:0] rf_14; // @[src/main/scala/nutcore/RF.scala 33:15]
  reg [63:0] rf_15; // @[src/main/scala/nutcore/RF.scala 33:15]
  reg [63:0] rf_16; // @[src/main/scala/nutcore/RF.scala 33:15]
  reg [63:0] rf_17; // @[src/main/scala/nutcore/RF.scala 33:15]
  reg [63:0] rf_18; // @[src/main/scala/nutcore/RF.scala 33:15]
  reg [63:0] rf_19; // @[src/main/scala/nutcore/RF.scala 33:15]
  reg [63:0] rf_20; // @[src/main/scala/nutcore/RF.scala 33:15]
  reg [63:0] rf_21; // @[src/main/scala/nutcore/RF.scala 33:15]
  reg [63:0] rf_22; // @[src/main/scala/nutcore/RF.scala 33:15]
  reg [63:0] rf_23; // @[src/main/scala/nutcore/RF.scala 33:15]
  reg [63:0] rf_24; // @[src/main/scala/nutcore/RF.scala 33:15]
  reg [63:0] rf_25; // @[src/main/scala/nutcore/RF.scala 33:15]
  reg [63:0] rf_26; // @[src/main/scala/nutcore/RF.scala 33:15]
  reg [63:0] rf_27; // @[src/main/scala/nutcore/RF.scala 33:15]
  reg [63:0] rf_28; // @[src/main/scala/nutcore/RF.scala 33:15]
  reg [63:0] rf_29; // @[src/main/scala/nutcore/RF.scala 33:15]
  reg [63:0] rf_30; // @[src/main/scala/nutcore/RF.scala 33:15]
  reg [63:0] rf_31; // @[src/main/scala/nutcore/RF.scala 33:15]
  wire  io_out_bits_data_src1_signBit = io_in_0_bits_cf_pc[38]; // @[src/main/scala/utils/BitUtils.scala 39:20]
  wire [24:0] _io_out_bits_data_src1_T_2 = io_out_bits_data_src1_signBit ? 25'h1ffffff : 25'h0; // @[src/main/scala/utils/BitUtils.scala 40:46]
  wire [63:0] _io_out_bits_data_src1_T_3 = {_io_out_bits_data_src1_T_2,io_in_0_bits_cf_pc}; // @[src/main/scala/utils/BitUtils.scala 40:41]
  wire  _io_out_bits_data_src1_T_4 = ~src1ForwardNextCycle; // @[src/main/scala/nutcore/backend/seq/ISU.scala 66:21]
  wire  _io_out_bits_data_src1_T_5 = src1Forward & ~src1ForwardNextCycle; // @[src/main/scala/nutcore/backend/seq/ISU.scala 66:18]
  wire  _io_out_bits_data_src1_T_10 = ~io_in_0_bits_ctrl_src1Type & _io_out_bits_data_src1_T_4 & ~src1Forward; // @[src/main/scala/nutcore/backend/seq/ISU.scala 67:76]
  wire [63:0] _GEN_1 = 5'h1 == io_in_0_bits_ctrl_rfSrc1 ? rf_1 : rf_0; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_2 = 5'h2 == io_in_0_bits_ctrl_rfSrc1 ? rf_2 : _GEN_1; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_3 = 5'h3 == io_in_0_bits_ctrl_rfSrc1 ? rf_3 : _GEN_2; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_4 = 5'h4 == io_in_0_bits_ctrl_rfSrc1 ? rf_4 : _GEN_3; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_5 = 5'h5 == io_in_0_bits_ctrl_rfSrc1 ? rf_5 : _GEN_4; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_6 = 5'h6 == io_in_0_bits_ctrl_rfSrc1 ? rf_6 : _GEN_5; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_7 = 5'h7 == io_in_0_bits_ctrl_rfSrc1 ? rf_7 : _GEN_6; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_8 = 5'h8 == io_in_0_bits_ctrl_rfSrc1 ? rf_8 : _GEN_7; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_9 = 5'h9 == io_in_0_bits_ctrl_rfSrc1 ? rf_9 : _GEN_8; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_10 = 5'ha == io_in_0_bits_ctrl_rfSrc1 ? rf_10 : _GEN_9; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_11 = 5'hb == io_in_0_bits_ctrl_rfSrc1 ? rf_11 : _GEN_10; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_12 = 5'hc == io_in_0_bits_ctrl_rfSrc1 ? rf_12 : _GEN_11; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_13 = 5'hd == io_in_0_bits_ctrl_rfSrc1 ? rf_13 : _GEN_12; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_14 = 5'he == io_in_0_bits_ctrl_rfSrc1 ? rf_14 : _GEN_13; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_15 = 5'hf == io_in_0_bits_ctrl_rfSrc1 ? rf_15 : _GEN_14; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_16 = 5'h10 == io_in_0_bits_ctrl_rfSrc1 ? rf_16 : _GEN_15; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_17 = 5'h11 == io_in_0_bits_ctrl_rfSrc1 ? rf_17 : _GEN_16; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_18 = 5'h12 == io_in_0_bits_ctrl_rfSrc1 ? rf_18 : _GEN_17; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_19 = 5'h13 == io_in_0_bits_ctrl_rfSrc1 ? rf_19 : _GEN_18; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_20 = 5'h14 == io_in_0_bits_ctrl_rfSrc1 ? rf_20 : _GEN_19; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_21 = 5'h15 == io_in_0_bits_ctrl_rfSrc1 ? rf_21 : _GEN_20; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_22 = 5'h16 == io_in_0_bits_ctrl_rfSrc1 ? rf_22 : _GEN_21; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_23 = 5'h17 == io_in_0_bits_ctrl_rfSrc1 ? rf_23 : _GEN_22; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_24 = 5'h18 == io_in_0_bits_ctrl_rfSrc1 ? rf_24 : _GEN_23; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_25 = 5'h19 == io_in_0_bits_ctrl_rfSrc1 ? rf_25 : _GEN_24; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_26 = 5'h1a == io_in_0_bits_ctrl_rfSrc1 ? rf_26 : _GEN_25; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_27 = 5'h1b == io_in_0_bits_ctrl_rfSrc1 ? rf_27 : _GEN_26; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_28 = 5'h1c == io_in_0_bits_ctrl_rfSrc1 ? rf_28 : _GEN_27; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_29 = 5'h1d == io_in_0_bits_ctrl_rfSrc1 ? rf_29 : _GEN_28; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_30 = 5'h1e == io_in_0_bits_ctrl_rfSrc1 ? rf_30 : _GEN_29; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_31 = 5'h1f == io_in_0_bits_ctrl_rfSrc1 ? rf_31 : _GEN_30; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _io_out_bits_data_src1_T_12 = io_in_0_bits_ctrl_rfSrc1 == 5'h0 ? 64'h0 : _GEN_31; // @[src/main/scala/nutcore/RF.scala 40:37]
  wire [63:0] _io_out_bits_data_src1_T_13 = io_in_0_bits_ctrl_src1Type ? _io_out_bits_data_src1_T_3 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src1_T_14 = src1ForwardNextCycle ? io_forward_wb_rfData : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src1_T_15 = _io_out_bits_data_src1_T_5 ? io_wb_rfData : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src1_T_16 = _io_out_bits_data_src1_T_10 ? _io_out_bits_data_src1_T_12 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src1_T_17 = _io_out_bits_data_src1_T_13 | _io_out_bits_data_src1_T_14; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src1_T_18 = _io_out_bits_data_src1_T_17 | _io_out_bits_data_src1_T_15; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_out_bits_data_src2_T_1 = ~src2ForwardNextCycle; // @[src/main/scala/nutcore/backend/seq/ISU.scala 72:21]
  wire  _io_out_bits_data_src2_T_2 = src2Forward & ~src2ForwardNextCycle; // @[src/main/scala/nutcore/backend/seq/ISU.scala 72:18]
  wire  _io_out_bits_data_src2_T_7 = ~io_in_0_bits_ctrl_src2Type & _io_out_bits_data_src2_T_1 & ~src2Forward; // @[src/main/scala/nutcore/backend/seq/ISU.scala 73:77]
  wire [63:0] _GEN_33 = 5'h1 == io_in_0_bits_ctrl_rfSrc2 ? rf_1 : rf_0; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_34 = 5'h2 == io_in_0_bits_ctrl_rfSrc2 ? rf_2 : _GEN_33; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_35 = 5'h3 == io_in_0_bits_ctrl_rfSrc2 ? rf_3 : _GEN_34; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_36 = 5'h4 == io_in_0_bits_ctrl_rfSrc2 ? rf_4 : _GEN_35; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_37 = 5'h5 == io_in_0_bits_ctrl_rfSrc2 ? rf_5 : _GEN_36; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_38 = 5'h6 == io_in_0_bits_ctrl_rfSrc2 ? rf_6 : _GEN_37; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_39 = 5'h7 == io_in_0_bits_ctrl_rfSrc2 ? rf_7 : _GEN_38; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_40 = 5'h8 == io_in_0_bits_ctrl_rfSrc2 ? rf_8 : _GEN_39; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_41 = 5'h9 == io_in_0_bits_ctrl_rfSrc2 ? rf_9 : _GEN_40; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_42 = 5'ha == io_in_0_bits_ctrl_rfSrc2 ? rf_10 : _GEN_41; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_43 = 5'hb == io_in_0_bits_ctrl_rfSrc2 ? rf_11 : _GEN_42; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_44 = 5'hc == io_in_0_bits_ctrl_rfSrc2 ? rf_12 : _GEN_43; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_45 = 5'hd == io_in_0_bits_ctrl_rfSrc2 ? rf_13 : _GEN_44; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_46 = 5'he == io_in_0_bits_ctrl_rfSrc2 ? rf_14 : _GEN_45; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_47 = 5'hf == io_in_0_bits_ctrl_rfSrc2 ? rf_15 : _GEN_46; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_48 = 5'h10 == io_in_0_bits_ctrl_rfSrc2 ? rf_16 : _GEN_47; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_49 = 5'h11 == io_in_0_bits_ctrl_rfSrc2 ? rf_17 : _GEN_48; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_50 = 5'h12 == io_in_0_bits_ctrl_rfSrc2 ? rf_18 : _GEN_49; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_51 = 5'h13 == io_in_0_bits_ctrl_rfSrc2 ? rf_19 : _GEN_50; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_52 = 5'h14 == io_in_0_bits_ctrl_rfSrc2 ? rf_20 : _GEN_51; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_53 = 5'h15 == io_in_0_bits_ctrl_rfSrc2 ? rf_21 : _GEN_52; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_54 = 5'h16 == io_in_0_bits_ctrl_rfSrc2 ? rf_22 : _GEN_53; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_55 = 5'h17 == io_in_0_bits_ctrl_rfSrc2 ? rf_23 : _GEN_54; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_56 = 5'h18 == io_in_0_bits_ctrl_rfSrc2 ? rf_24 : _GEN_55; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_57 = 5'h19 == io_in_0_bits_ctrl_rfSrc2 ? rf_25 : _GEN_56; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_58 = 5'h1a == io_in_0_bits_ctrl_rfSrc2 ? rf_26 : _GEN_57; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_59 = 5'h1b == io_in_0_bits_ctrl_rfSrc2 ? rf_27 : _GEN_58; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_60 = 5'h1c == io_in_0_bits_ctrl_rfSrc2 ? rf_28 : _GEN_59; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_61 = 5'h1d == io_in_0_bits_ctrl_rfSrc2 ? rf_29 : _GEN_60; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_62 = 5'h1e == io_in_0_bits_ctrl_rfSrc2 ? rf_30 : _GEN_61; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _GEN_63 = 5'h1f == io_in_0_bits_ctrl_rfSrc2 ? rf_31 : _GEN_62; // @[src/main/scala/nutcore/RF.scala 40:{37,37}]
  wire [63:0] _io_out_bits_data_src2_T_9 = io_in_0_bits_ctrl_rfSrc2 == 5'h0 ? 64'h0 : _GEN_63; // @[src/main/scala/nutcore/RF.scala 40:37]
  wire [63:0] _io_out_bits_data_src2_T_10 = io_in_0_bits_ctrl_src2Type ? io_in_0_bits_data_imm : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src2_T_11 = src2ForwardNextCycle ? io_forward_wb_rfData : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src2_T_12 = _io_out_bits_data_src2_T_2 ? io_wb_rfData : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src2_T_13 = _io_out_bits_data_src2_T_7 ? _io_out_bits_data_src2_T_9 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src2_T_14 = _io_out_bits_data_src2_T_10 | _io_out_bits_data_src2_T_11; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src2_T_15 = _io_out_bits_data_src2_T_14 | _io_out_bits_data_src2_T_12; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _T = io_wb_rfDest != 5'h0; // @[src/main/scala/nutcore/RF.scala 42:15]
  wire  _wbClearMask_T_3 = _T & io_wb_rfDest == io_forward_wb_rfDest & forwardRfWen; // @[src/main/scala/nutcore/backend/seq/ISU.scala 41:100]
  wire [62:0] _wbClearMask_T_6 = 63'h1 << io_wb_rfDest; // @[src/main/scala/nutcore/RF.scala 52:39]
  wire [31:0] wbClearMask = io_wb_rfWen & ~_wbClearMask_T_3 ? _wbClearMask_T_6[31:0] : 32'h0; // @[src/main/scala/nutcore/backend/seq/ISU.scala 85:24]
  wire  _isuFireSetMask_T = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [62:0] _isuFireSetMask_T_1 = 63'h1 << io_in_0_bits_ctrl_rfDest; // @[src/main/scala/nutcore/RF.scala 52:39]
  wire [31:0] isuFireSetMask = _isuFireSetMask_T ? _isuFireSetMask_T_1[31:0] : 32'h0; // @[src/main/scala/nutcore/backend/seq/ISU.scala 87:27]
  wire [31:0] _busy_T_5 = ~wbClearMask; // @[src/main/scala/nutcore/RF.scala 58:26]
  wire [31:0] _busy_T_6 = busy & _busy_T_5; // @[src/main/scala/nutcore/RF.scala 58:24]
  wire [31:0] _busy_T_7 = _busy_T_6 | isuFireSetMask; // @[src/main/scala/nutcore/RF.scala 58:38]
  wire [31:0] _busy_T_9 = {_busy_T_7[31:1],1'h0}; // @[src/main/scala/nutcore/RF.scala 58:16]
  wire  _T_9 = io_in_0_valid & ~io_out_valid; // @[src/main/scala/nutcore/backend/seq/ISU.scala 97:40]
  wire  _T_12 = io_out_valid & ~_isuFireSetMask_T; // @[src/main/scala/nutcore/backend/seq/ISU.scala 98:38]
  wire  _T_13 = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  assign io_in_0_ready = ~io_in_0_valid | _isuFireSetMask_T; // @[src/main/scala/nutcore/backend/seq/ISU.scala 91:37]
  assign io_out_valid = io_in_0_valid & src1Ready & src2Ready; // @[src/main/scala/nutcore/backend/seq/ISU.scala 58:47]
  assign io_out_bits_cf_instr = io_in_0_bits_cf_instr; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_pc = io_in_0_bits_cf_pc; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_pnpc = io_in_0_bits_cf_pnpc; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_exceptionVec_1 = io_in_0_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_exceptionVec_2 = io_in_0_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_0 = io_in_0_bits_cf_intrVec_0; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_1 = io_in_0_bits_cf_intrVec_1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_2 = io_in_0_bits_cf_intrVec_2; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_3 = io_in_0_bits_cf_intrVec_3; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_4 = io_in_0_bits_cf_intrVec_4; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_5 = io_in_0_bits_cf_intrVec_5; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_6 = io_in_0_bits_cf_intrVec_6; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_7 = io_in_0_bits_cf_intrVec_7; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_8 = io_in_0_bits_cf_intrVec_8; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_9 = io_in_0_bits_cf_intrVec_9; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_10 = io_in_0_bits_cf_intrVec_10; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_11 = io_in_0_bits_cf_intrVec_11; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_brIdx = io_in_0_bits_cf_brIdx; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_ctrl_fuType = io_in_0_bits_ctrl_fuType; // @[src/main/scala/nutcore/backend/seq/ISU.scala 78:20]
  assign io_out_bits_ctrl_fuOpType = io_in_0_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/seq/ISU.scala 78:20]
  assign io_out_bits_ctrl_rfSrc1 = io_in_0_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 78:20]
  assign io_out_bits_ctrl_rfSrc2 = io_in_0_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/backend/seq/ISU.scala 78:20]
  assign io_out_bits_ctrl_rfWen = io_in_0_bits_ctrl_rfWen; // @[src/main/scala/nutcore/backend/seq/ISU.scala 78:20]
  assign io_out_bits_ctrl_rfDest = io_in_0_bits_ctrl_rfDest; // @[src/main/scala/nutcore/backend/seq/ISU.scala 78:20]
  assign io_out_bits_data_src1 = _io_out_bits_data_src1_T_18 | _io_out_bits_data_src1_T_16; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_out_bits_data_src2 = _io_out_bits_data_src2_T_15 | _io_out_bits_data_src2_T_13; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_out_bits_data_imm = io_in_0_bits_data_imm; // @[src/main/scala/nutcore/backend/seq/ISU.scala 75:25]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 50:21]
      busy <= 32'h0; // @[src/main/scala/nutcore/RF.scala 50:21]
    end else if (io_flush) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 88:19]
      busy <= 32'h0; // @[src/main/scala/nutcore/RF.scala 58:10]
    end else begin
      busy <= _busy_T_9; // @[src/main/scala/nutcore/RF.scala 58:10]
    end
    if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (io_wb_rfDest != 5'h0) begin // @[src/main/scala/nutcore/RF.scala 42:23]
        if (5'h0 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 43:16]
          rf_0 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 43:16]
        end else begin
          rf_0 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 35:9]
        end
      end else begin
        rf_0 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 35:9]
      end
    end else begin
      rf_0 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 35:9]
    end
    if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (io_wb_rfDest != 5'h0) begin // @[src/main/scala/nutcore/RF.scala 42:23]
        if (5'h1 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 43:16]
          rf_1 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 43:16]
        end
      end
    end
    if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (io_wb_rfDest != 5'h0) begin // @[src/main/scala/nutcore/RF.scala 42:23]
        if (5'h2 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 43:16]
          rf_2 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 43:16]
        end
      end
    end
    if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (io_wb_rfDest != 5'h0) begin // @[src/main/scala/nutcore/RF.scala 42:23]
        if (5'h3 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 43:16]
          rf_3 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 43:16]
        end
      end
    end
    if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (io_wb_rfDest != 5'h0) begin // @[src/main/scala/nutcore/RF.scala 42:23]
        if (5'h4 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 43:16]
          rf_4 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 43:16]
        end
      end
    end
    if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (io_wb_rfDest != 5'h0) begin // @[src/main/scala/nutcore/RF.scala 42:23]
        if (5'h5 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 43:16]
          rf_5 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 43:16]
        end
      end
    end
    if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (io_wb_rfDest != 5'h0) begin // @[src/main/scala/nutcore/RF.scala 42:23]
        if (5'h6 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 43:16]
          rf_6 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 43:16]
        end
      end
    end
    if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (io_wb_rfDest != 5'h0) begin // @[src/main/scala/nutcore/RF.scala 42:23]
        if (5'h7 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 43:16]
          rf_7 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 43:16]
        end
      end
    end
    if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (io_wb_rfDest != 5'h0) begin // @[src/main/scala/nutcore/RF.scala 42:23]
        if (5'h8 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 43:16]
          rf_8 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 43:16]
        end
      end
    end
    if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (io_wb_rfDest != 5'h0) begin // @[src/main/scala/nutcore/RF.scala 42:23]
        if (5'h9 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 43:16]
          rf_9 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 43:16]
        end
      end
    end
    if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (io_wb_rfDest != 5'h0) begin // @[src/main/scala/nutcore/RF.scala 42:23]
        if (5'ha == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 43:16]
          rf_10 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 43:16]
        end
      end
    end
    if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (io_wb_rfDest != 5'h0) begin // @[src/main/scala/nutcore/RF.scala 42:23]
        if (5'hb == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 43:16]
          rf_11 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 43:16]
        end
      end
    end
    if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (io_wb_rfDest != 5'h0) begin // @[src/main/scala/nutcore/RF.scala 42:23]
        if (5'hc == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 43:16]
          rf_12 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 43:16]
        end
      end
    end
    if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (io_wb_rfDest != 5'h0) begin // @[src/main/scala/nutcore/RF.scala 42:23]
        if (5'hd == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 43:16]
          rf_13 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 43:16]
        end
      end
    end
    if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (io_wb_rfDest != 5'h0) begin // @[src/main/scala/nutcore/RF.scala 42:23]
        if (5'he == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 43:16]
          rf_14 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 43:16]
        end
      end
    end
    if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (io_wb_rfDest != 5'h0) begin // @[src/main/scala/nutcore/RF.scala 42:23]
        if (5'hf == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 43:16]
          rf_15 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 43:16]
        end
      end
    end
    if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (io_wb_rfDest != 5'h0) begin // @[src/main/scala/nutcore/RF.scala 42:23]
        if (5'h10 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 43:16]
          rf_16 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 43:16]
        end
      end
    end
    if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (io_wb_rfDest != 5'h0) begin // @[src/main/scala/nutcore/RF.scala 42:23]
        if (5'h11 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 43:16]
          rf_17 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 43:16]
        end
      end
    end
    if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (io_wb_rfDest != 5'h0) begin // @[src/main/scala/nutcore/RF.scala 42:23]
        if (5'h12 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 43:16]
          rf_18 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 43:16]
        end
      end
    end
    if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (io_wb_rfDest != 5'h0) begin // @[src/main/scala/nutcore/RF.scala 42:23]
        if (5'h13 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 43:16]
          rf_19 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 43:16]
        end
      end
    end
    if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (io_wb_rfDest != 5'h0) begin // @[src/main/scala/nutcore/RF.scala 42:23]
        if (5'h14 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 43:16]
          rf_20 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 43:16]
        end
      end
    end
    if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (io_wb_rfDest != 5'h0) begin // @[src/main/scala/nutcore/RF.scala 42:23]
        if (5'h15 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 43:16]
          rf_21 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 43:16]
        end
      end
    end
    if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (io_wb_rfDest != 5'h0) begin // @[src/main/scala/nutcore/RF.scala 42:23]
        if (5'h16 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 43:16]
          rf_22 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 43:16]
        end
      end
    end
    if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (io_wb_rfDest != 5'h0) begin // @[src/main/scala/nutcore/RF.scala 42:23]
        if (5'h17 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 43:16]
          rf_23 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 43:16]
        end
      end
    end
    if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (io_wb_rfDest != 5'h0) begin // @[src/main/scala/nutcore/RF.scala 42:23]
        if (5'h18 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 43:16]
          rf_24 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 43:16]
        end
      end
    end
    if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (io_wb_rfDest != 5'h0) begin // @[src/main/scala/nutcore/RF.scala 42:23]
        if (5'h19 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 43:16]
          rf_25 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 43:16]
        end
      end
    end
    if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (io_wb_rfDest != 5'h0) begin // @[src/main/scala/nutcore/RF.scala 42:23]
        if (5'h1a == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 43:16]
          rf_26 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 43:16]
        end
      end
    end
    if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (io_wb_rfDest != 5'h0) begin // @[src/main/scala/nutcore/RF.scala 42:23]
        if (5'h1b == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 43:16]
          rf_27 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 43:16]
        end
      end
    end
    if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (io_wb_rfDest != 5'h0) begin // @[src/main/scala/nutcore/RF.scala 42:23]
        if (5'h1c == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 43:16]
          rf_28 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 43:16]
        end
      end
    end
    if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (io_wb_rfDest != 5'h0) begin // @[src/main/scala/nutcore/RF.scala 42:23]
        if (5'h1d == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 43:16]
          rf_29 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 43:16]
        end
      end
    end
    if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (io_wb_rfDest != 5'h0) begin // @[src/main/scala/nutcore/RF.scala 42:23]
        if (5'h1e == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 43:16]
          rf_30 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 43:16]
        end
      end
    end
    if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (io_wb_rfDest != 5'h0) begin // @[src/main/scala/nutcore/RF.scala 42:23]
        if (5'h1f == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 43:16]
          rf_31 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 43:16]
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  busy = _RAND_0[31:0];
  _RAND_1 = {2{`RANDOM}};
  rf_0 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  rf_1 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  rf_2 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  rf_3 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  rf_4 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  rf_5 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  rf_6 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  rf_7 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  rf_8 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  rf_9 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  rf_10 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  rf_11 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  rf_12 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  rf_13 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  rf_14 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  rf_15 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  rf_16 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  rf_17 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  rf_18 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  rf_19 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  rf_20 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  rf_21 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  rf_22 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  rf_23 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  rf_24 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  rf_25 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  rf_26 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  rf_27 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  rf_28 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  rf_29 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  rf_30 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  rf_31 = _RAND_32[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ALU(
  input         clock,
  input         reset,
  input         io_in_valid, // @[src/main/scala/nutcore/backend/fu/ALU.scala 76:14]
  input  [63:0] io_in_bits_src1, // @[src/main/scala/nutcore/backend/fu/ALU.scala 76:14]
  input  [63:0] io_in_bits_src2, // @[src/main/scala/nutcore/backend/fu/ALU.scala 76:14]
  input  [6:0]  io_in_bits_func, // @[src/main/scala/nutcore/backend/fu/ALU.scala 76:14]
  input         io_out_ready, // @[src/main/scala/nutcore/backend/fu/ALU.scala 76:14]
  output        io_out_valid, // @[src/main/scala/nutcore/backend/fu/ALU.scala 76:14]
  output [63:0] io_out_bits, // @[src/main/scala/nutcore/backend/fu/ALU.scala 76:14]
  input  [63:0] io_cfIn_instr, // @[src/main/scala/nutcore/backend/fu/ALU.scala 76:14]
  input  [38:0] io_cfIn_pc, // @[src/main/scala/nutcore/backend/fu/ALU.scala 76:14]
  input  [38:0] io_cfIn_pnpc, // @[src/main/scala/nutcore/backend/fu/ALU.scala 76:14]
  input  [3:0]  io_cfIn_brIdx, // @[src/main/scala/nutcore/backend/fu/ALU.scala 76:14]
  output [38:0] io_redirect_target, // @[src/main/scala/nutcore/backend/fu/ALU.scala 76:14]
  output        io_redirect_valid, // @[src/main/scala/nutcore/backend/fu/ALU.scala 76:14]
  input  [63:0] io_offset, // @[src/main/scala/nutcore/backend/fu/ALU.scala 76:14]
  output        _T_2_0,
  output        REG_0_valid,
  output [38:0] REG_0_pc,
  output        REG_0_isMissPredict,
  output [38:0] REG_0_actualTarget,
  output        REG_0_actualTaken,
  output [6:0]  REG_0_fuOpType,
  output [1:0]  REG_0_btbType,
  output        REG_0_isRVC
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  isAdderSub = ~io_in_bits_func[6]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 87:20]
  wire [63:0] _adderRes_T_1 = isAdderSub ? 64'hffffffffffffffff : 64'h0; // @[src/main/scala/nutcore/backend/fu/ALU.scala 88:39]
  wire [63:0] _adderRes_T_2 = io_in_bits_src2 ^ _adderRes_T_1; // @[src/main/scala/nutcore/backend/fu/ALU.scala 88:33]
  wire [64:0] _adderRes_T_3 = io_in_bits_src1 + _adderRes_T_2; // @[src/main/scala/nutcore/backend/fu/ALU.scala 88:24]
  wire [64:0] _GEN_0 = {{64'd0}, isAdderSub}; // @[src/main/scala/nutcore/backend/fu/ALU.scala 88:60]
  wire [64:0] adderRes = _adderRes_T_3 + _GEN_0; // @[src/main/scala/nutcore/backend/fu/ALU.scala 88:60]
  wire [63:0] xorRes = io_in_bits_src1 ^ io_in_bits_src2; // @[src/main/scala/nutcore/backend/fu/ALU.scala 89:21]
  wire  sltu = ~adderRes[64]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 90:14]
  wire  slt = xorRes[63] ^ sltu; // @[src/main/scala/nutcore/backend/fu/ALU.scala 91:28]
  wire [63:0] _shsrc1_T_2 = {32'h0,io_in_bits_src1[31:0]}; // @[src/main/scala/utils/BitUtils.scala 47:41]
  wire  shsrc1_signBit = io_in_bits_src1[31]; // @[src/main/scala/utils/BitUtils.scala 39:20]
  wire [31:0] _shsrc1_T_5 = shsrc1_signBit ? 32'hffffffff : 32'h0; // @[src/main/scala/utils/BitUtils.scala 40:46]
  wire [63:0] _shsrc1_T_6 = {_shsrc1_T_5,io_in_bits_src1[31:0]}; // @[src/main/scala/utils/BitUtils.scala 40:41]
  wire [63:0] _shsrc1_T_8 = 7'h25 == io_in_bits_func ? _shsrc1_T_2 : io_in_bits_src1; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [63:0] shsrc1 = 7'h2d == io_in_bits_func ? _shsrc1_T_6 : _shsrc1_T_8; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [5:0] shamt = io_in_bits_func[5] ? {{1'd0}, io_in_bits_src2[4:0]} : io_in_bits_src2[5:0]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 97:18]
  wire [126:0] _GEN_4 = {{63'd0}, shsrc1}; // @[src/main/scala/nutcore/backend/fu/ALU.scala 99:33]
  wire [126:0] _res_T_1 = _GEN_4 << shamt; // @[src/main/scala/nutcore/backend/fu/ALU.scala 99:33]
  wire [63:0] _res_T_3 = {63'h0,slt}; // @[src/main/scala/utils/BitUtils.scala 47:41]
  wire [63:0] _res_T_4 = {63'h0,sltu}; // @[src/main/scala/utils/BitUtils.scala 47:41]
  wire [63:0] _res_T_5 = shsrc1 >> shamt; // @[src/main/scala/nutcore/backend/fu/ALU.scala 103:32]
  wire [63:0] _res_T_6 = io_in_bits_src1 | io_in_bits_src2; // @[src/main/scala/nutcore/backend/fu/ALU.scala 104:30]
  wire [63:0] _res_T_7 = io_in_bits_src1 & io_in_bits_src2; // @[src/main/scala/nutcore/backend/fu/ALU.scala 105:30]
  wire [63:0] _res_T_8 = 7'h2d == io_in_bits_func ? _shsrc1_T_6 : _shsrc1_T_8; // @[src/main/scala/nutcore/backend/fu/ALU.scala 106:32]
  wire [63:0] _res_T_10 = $signed(_res_T_8) >>> shamt; // @[src/main/scala/nutcore/backend/fu/ALU.scala 106:49]
  wire [63:0] _res_T_12 = io_in_bits_src1 - io_in_bits_src2; // @[src/main/scala/nutcore/backend/fu/ALU.scala 107:45]
  wire [63:0] _res_T_14 = {1'h0,_res_T_12[62:0]}; // @[src/main/scala/nutcore/backend/fu/ALU.scala 107:27]
  wire [64:0] _res_T_16 = 4'h1 == io_in_bits_func[3:0] ? {{1'd0}, _res_T_1[63:0]} : adderRes; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_18 = 4'h2 == io_in_bits_func[3:0] ? {{1'd0}, _res_T_3} : _res_T_16; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_20 = 4'h3 == io_in_bits_func[3:0] ? {{1'd0}, _res_T_4} : _res_T_18; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_22 = 4'h4 == io_in_bits_func[3:0] ? {{1'd0}, xorRes} : _res_T_20; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_24 = 4'h5 == io_in_bits_func[3:0] ? {{1'd0}, _res_T_5} : _res_T_22; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_26 = 4'h6 == io_in_bits_func[3:0] ? {{1'd0}, _res_T_6} : _res_T_24; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_28 = 4'h7 == io_in_bits_func[3:0] ? {{1'd0}, _res_T_7} : _res_T_26; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_30 = 4'hd == io_in_bits_func[3:0] ? {{1'd0}, _res_T_10} : _res_T_28; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] res = 4'hb == io_in_bits_func[3:0] ? {{1'd0}, _res_T_14} : _res_T_30; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  aluRes_signBit = res[31]; // @[src/main/scala/utils/BitUtils.scala 39:20]
  wire [31:0] _aluRes_T_3 = aluRes_signBit ? 32'hffffffff : 32'h0; // @[src/main/scala/utils/BitUtils.scala 40:46]
  wire [63:0] _aluRes_T_4 = {_aluRes_T_3,res[31:0]}; // @[src/main/scala/utils/BitUtils.scala 40:41]
  wire [64:0] aluRes = io_in_bits_func[5] ? {{1'd0}, _aluRes_T_4} : res; // @[src/main/scala/nutcore/backend/fu/ALU.scala 109:19]
  wire  _T_1 = ~(|xorRes); // @[src/main/scala/nutcore/backend/fu/ALU.scala 112:48]
  wire  isBranch = ~io_in_bits_func[3]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 63:30]
  wire  isBru = io_in_bits_func[4]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 62:31]
  wire  _taken_T_1 = 2'h0 == io_in_bits_func[2:1]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _taken_T_2 = 2'h2 == io_in_bits_func[2:1]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _taken_T_3 = 2'h3 == io_in_bits_func[2:1]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _taken_T_8 = _taken_T_1 & _T_1 | _taken_T_2 & slt | _taken_T_3 & sltu; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  taken = _taken_T_8 ^ io_in_bits_func[0]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 119:72]
  wire [63:0] _GEN_1 = {{25'd0}, io_cfIn_pc}; // @[src/main/scala/nutcore/backend/fu/ALU.scala 120:41]
  wire [63:0] _target_T_1 = _GEN_1 + io_offset; // @[src/main/scala/nutcore/backend/fu/ALU.scala 120:41]
  wire [64:0] _target_T_2 = isBranch ? {{1'd0}, _target_T_1} : adderRes; // @[src/main/scala/nutcore/backend/fu/ALU.scala 120:19]
  wire [38:0] target = _target_T_2[38:0]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 120:63]
  wire  _targetAssume_T_3 = target[1:0] == 2'h0; // @[src/main/scala/nutcore/backend/fu/ALU.scala 121:59]
  wire  targetAssume = ~(isBranch & taken) | target[1:0] == 2'h0; // @[src/main/scala/nutcore/backend/fu/ALU.scala 121:43]
  wire  _jumpAssume_T_4 = isBru & ~isBranch; // @[src/main/scala/nutcore/backend/fu/ALU.scala 64:40]
  wire  jumpAssume = ~_jumpAssume_T_4 | _targetAssume_T_3; // @[src/main/scala/nutcore/backend/fu/ALU.scala 122:46]
  wire  _T_2 = targetAssume & jumpAssume; // @[src/main/scala/nutcore/backend/fu/ALU.scala 124:38]
  wire  _predictWrong_T_1 = ~taken & isBranch; // @[src/main/scala/nutcore/backend/fu/ALU.scala 131:33]
  wire  predictWrong = ~taken & isBranch ? io_cfIn_brIdx[0] : ~io_cfIn_brIdx[0] | io_redirect_target != io_cfIn_pnpc; // @[src/main/scala/nutcore/backend/fu/ALU.scala 131:25]
  wire  isRVC = io_cfIn_instr[1:0] != 2'h3; // @[src/main/scala/nutcore/backend/fu/ALU.scala 132:35]
  wire  _T_13 = ~isRVC; // @[src/main/scala/nutcore/backend/fu/ALU.scala 134:55]
  wire [38:0] _io_redirect_target_T_3 = io_cfIn_pc + 39'h2; // @[src/main/scala/nutcore/backend/fu/ALU.scala 135:71]
  wire [38:0] _io_redirect_target_T_5 = io_cfIn_pc + 39'h4; // @[src/main/scala/nutcore/backend/fu/ALU.scala 135:89]
  wire [38:0] _io_redirect_target_T_6 = isRVC ? _io_redirect_target_T_3 : _io_redirect_target_T_5; // @[src/main/scala/nutcore/backend/fu/ALU.scala 135:52]
  wire  _io_redirect_valid_T = io_in_valid & isBru; // @[src/main/scala/nutcore/backend/fu/ALU.scala 137:30]
  wire  _io_redirect_valid_T_1 = io_in_valid & isBru & predictWrong; // @[src/main/scala/nutcore/backend/fu/ALU.scala 137:39]
  wire  io_out_bits_signBit = io_cfIn_pc[38]; // @[src/main/scala/utils/BitUtils.scala 39:20]
  wire [24:0] _io_out_bits_T_2 = io_out_bits_signBit ? 25'h1ffffff : 25'h0; // @[src/main/scala/utils/BitUtils.scala 40:46]
  wire [63:0] _io_out_bits_T_3 = {_io_out_bits_T_2,io_cfIn_pc}; // @[src/main/scala/utils/BitUtils.scala 40:41]
  wire [63:0] _io_out_bits_T_5 = _io_out_bits_T_3 + 64'h4; // @[src/main/scala/nutcore/backend/fu/ALU.scala 143:71]
  wire [63:0] _io_out_bits_T_10 = _io_out_bits_T_3 + 64'h2; // @[src/main/scala/nutcore/backend/fu/ALU.scala 143:108]
  wire [63:0] _io_out_bits_T_11 = _T_13 ? _io_out_bits_T_5 : _io_out_bits_T_10; // @[src/main/scala/nutcore/backend/fu/ALU.scala 143:32]
  wire [64:0] _io_out_bits_T_12 = isBru ? {{1'd0}, _io_out_bits_T_11} : aluRes; // @[src/main/scala/nutcore/backend/fu/ALU.scala 143:21]
  wire  _T_36 = io_in_bits_func == 7'h58 | io_in_bits_func == 7'h5c; // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:180]
  wire  _T_37 = io_in_bits_func == 7'h5a; // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:214]
  wire  _T_38 = io_in_bits_func == 7'h5e; // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:239]
  wire  _T_57 = 7'h5c == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _T_58 = 7'h5e == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _T_59 = 7'h58 == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _T_60 = 7'h5a == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [1:0] _T_68 = _T_58 ? 2'h3 : 2'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _T_70 = _T_60 ? 2'h2 : 2'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _GEN_2 = {{1'd0}, _T_57}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _T_77 = _GEN_2 | _T_68; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _GEN_3 = {{1'd0}, _T_59}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _T_78 = _T_77 | _GEN_3; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  reg  REG_valid; // @[src/main/scala/nutcore/backend/fu/ALU.scala 170:34]
  reg [38:0] REG_pc; // @[src/main/scala/nutcore/backend/fu/ALU.scala 170:34]
  reg  REG_isMissPredict; // @[src/main/scala/nutcore/backend/fu/ALU.scala 170:34]
  reg [38:0] REG_actualTarget; // @[src/main/scala/nutcore/backend/fu/ALU.scala 170:34]
  reg  REG_actualTaken; // @[src/main/scala/nutcore/backend/fu/ALU.scala 170:34]
  reg [6:0] REG_fuOpType; // @[src/main/scala/nutcore/backend/fu/ALU.scala 170:34]
  reg [1:0] REG_btbType; // @[src/main/scala/nutcore/backend/fu/ALU.scala 170:34]
  reg  REG_isRVC; // @[src/main/scala/nutcore/backend/fu/ALU.scala 170:34]
  wire  right = _io_redirect_valid_T & ~predictWrong; // @[src/main/scala/nutcore/backend/fu/ALU.scala 172:32]
  wire  _T_85 = right & isBranch; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:33]
  wire  _T_86 = _io_redirect_valid_T_1 & isBranch; // @[src/main/scala/nutcore/backend/fu/ALU.scala 175:33]
  wire  _T_90 = _T_86 & io_cfIn_pc[2:0] == 3'h0; // @[src/main/scala/nutcore/backend/fu/ALU.scala 176:45]
  wire  _T_91 = _T_86 & io_cfIn_pc[2:0] == 3'h0 & isRVC; // @[src/main/scala/nutcore/backend/fu/ALU.scala 176:73]
  wire  _T_97 = _T_90 & _T_13; // @[src/main/scala/nutcore/backend/fu/ALU.scala 177:73]
  wire  _T_101 = _T_86 & io_cfIn_pc[2:0] == 3'h2; // @[src/main/scala/nutcore/backend/fu/ALU.scala 178:45]
  wire  _T_102 = _T_86 & io_cfIn_pc[2:0] == 3'h2 & isRVC; // @[src/main/scala/nutcore/backend/fu/ALU.scala 178:73]
  wire  _T_108 = _T_101 & _T_13; // @[src/main/scala/nutcore/backend/fu/ALU.scala 179:73]
  wire  _T_112 = _T_86 & io_cfIn_pc[2:0] == 3'h4; // @[src/main/scala/nutcore/backend/fu/ALU.scala 180:45]
  wire  _T_113 = _T_86 & io_cfIn_pc[2:0] == 3'h4 & isRVC; // @[src/main/scala/nutcore/backend/fu/ALU.scala 180:73]
  wire  _T_119 = _T_112 & _T_13; // @[src/main/scala/nutcore/backend/fu/ALU.scala 181:73]
  wire  _T_123 = _T_86 & io_cfIn_pc[2:0] == 3'h6; // @[src/main/scala/nutcore/backend/fu/ALU.scala 182:45]
  wire  _T_124 = _T_86 & io_cfIn_pc[2:0] == 3'h6 & isRVC; // @[src/main/scala/nutcore/backend/fu/ALU.scala 182:73]
  wire  _T_130 = _T_123 & _T_13; // @[src/main/scala/nutcore/backend/fu/ALU.scala 183:73]
  wire  _T_134 = right & _T_36; // @[src/main/scala/nutcore/backend/fu/ALU.scala 184:33]
  wire  _T_138 = _io_redirect_valid_T_1 & _T_36; // @[src/main/scala/nutcore/backend/fu/ALU.scala 185:33]
  wire  _T_140 = right & _T_37; // @[src/main/scala/nutcore/backend/fu/ALU.scala 186:33]
  wire  _T_142 = _io_redirect_valid_T_1 & _T_37; // @[src/main/scala/nutcore/backend/fu/ALU.scala 187:33]
  wire  _T_144 = right & _T_38; // @[src/main/scala/nutcore/backend/fu/ALU.scala 188:33]
  wire  _T_146 = _io_redirect_valid_T_1 & _T_38; // @[src/main/scala/nutcore/backend/fu/ALU.scala 189:33]
  assign io_out_valid = io_in_valid; // @[src/main/scala/nutcore/backend/fu/ALU.scala 157:16]
  assign io_out_bits = _io_out_bits_T_12[63:0]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 143:15]
  assign io_redirect_target = _predictWrong_T_1 ? _io_redirect_target_T_6 : target; // @[src/main/scala/nutcore/backend/fu/ALU.scala 135:28]
  assign io_redirect_valid = io_in_valid & isBru & predictWrong; // @[src/main/scala/nutcore/backend/fu/ALU.scala 137:39]
  assign _T_2_0 = _T_2;
  assign REG_0_valid = REG_valid;
  assign REG_0_pc = REG_pc;
  assign REG_0_isMissPredict = REG_isMissPredict;
  assign REG_0_actualTarget = REG_actualTarget;
  assign REG_0_actualTaken = REG_actualTaken;
  assign REG_0_fuOpType = REG_fuOpType;
  assign REG_0_btbType = REG_btbType;
  assign REG_0_isRVC = REG_isRVC;
  always @(posedge clock) begin
    REG_valid <= io_in_valid & isBru; // @[src/main/scala/nutcore/backend/fu/ALU.scala 160:31]
    REG_pc <= io_cfIn_pc; // @[src/main/scala/nutcore/backend/fu/ALU.scala 159:30 161:19]
    if (~taken & isBranch) begin // @[src/main/scala/nutcore/backend/fu/ALU.scala 131:25]
      REG_isMissPredict <= io_cfIn_brIdx[0];
    end else begin
      REG_isMissPredict <= ~io_cfIn_brIdx[0] | io_redirect_target != io_cfIn_pnpc;
    end
    REG_actualTarget <= _target_T_2[38:0]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 120:63]
    REG_actualTaken <= _taken_T_8 ^ io_in_bits_func[0]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 119:72]
    REG_fuOpType <= io_in_bits_func; // @[src/main/scala/nutcore/backend/fu/ALU.scala 159:30 165:25]
    REG_btbType <= _T_78 | _T_70; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
    REG_isRVC <= io_cfIn_instr[1:0] != 2'h3; // @[src/main/scala/nutcore/backend/fu/ALU.scala 132:35]
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_cfIn_instr[1:0] == 2'h3 | isRVC | ~io_in_valid)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ALU.scala:133 assert(io.cfIn.instr(1,0) === \"b11\".U || isRVC || !valid)\n"); // @[src/main/scala/nutcore/backend/fu/ALU.scala 133:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG_valid = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  REG_pc = _RAND_1[38:0];
  _RAND_2 = {1{`RANDOM}};
  REG_isMissPredict = _RAND_2[0:0];
  _RAND_3 = {2{`RANDOM}};
  REG_actualTarget = _RAND_3[38:0];
  _RAND_4 = {1{`RANDOM}};
  REG_actualTaken = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  REG_fuOpType = _RAND_5[6:0];
  _RAND_6 = {1{`RANDOM}};
  REG_btbType = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  REG_isRVC = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(io_cfIn_instr[1:0] == 2'h3 | isRVC | ~io_in_valid); // @[src/main/scala/nutcore/backend/fu/ALU.scala 133:9]
    end
  end
endmodule
module LSExecUnit(
  input         clock,
  input         reset,
  input         io__in_valid, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 290:14]
  input  [63:0] io__in_bits_src1, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 290:14]
  input  [6:0]  io__in_bits_func, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 290:14]
  input         io__out_ready, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 290:14]
  output        io__out_valid, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 290:14]
  output [63:0] io__out_bits, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 290:14]
  input  [63:0] io__wdata, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 290:14]
  input         io__dmem_req_ready, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 290:14]
  output        io__dmem_req_valid, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 290:14]
  output [38:0] io__dmem_req_bits_addr, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 290:14]
  output [2:0]  io__dmem_req_bits_size, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 290:14]
  output [3:0]  io__dmem_req_bits_cmd, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 290:14]
  output [7:0]  io__dmem_req_bits_wmask, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 290:14]
  output [63:0] io__dmem_req_bits_wdata, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 290:14]
  output        io__dmem_resp_ready, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 290:14]
  input         io__dmem_resp_valid, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 290:14]
  input  [63:0] io__dmem_resp_bits_rdata, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 290:14]
  output        io__isMMIO, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 290:14]
  output        io__loadAddrMisaligned, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 290:14]
  output        io__storeAddrMisaligned, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 290:14]
  input         ISAMO2,
  output [63:0] io_in_bits_src1
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] addrLatch; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 333:26]
  wire  isStore = io__in_valid & io__in_bits_func[3]; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 334:23]
  wire  _partialLoad_T = ~isStore; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 335:21]
  wire  partialLoad = ~isStore & io__in_bits_func != 7'h3; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 335:30]
  reg [1:0] state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 338:22]
  wire  _T_6 = io__dmem_req_ready & io__dmem_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _T_16 = io__dmem_resp_ready & io__dmem_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [1:0] _state_T = partialLoad ? 2'h3 : 2'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 361:60]
  wire [1:0] _GEN_4 = _T_16 ? _state_T : state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 338:22 361:{46,54}]
  wire [1:0] _GEN_5 = 2'h3 == state ? 2'h0 : state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 351:18 338:22 362:32]
  wire [63:0] _reqWdata_T_3 = {io__wdata[7:0],io__wdata[7:0],io__wdata[7:0],io__wdata[7:0],io__wdata[7:0],io__wdata[7:0]
    ,io__wdata[7:0],io__wdata[7:0]}; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 310:22]
  wire [63:0] _reqWdata_T_6 = {io__wdata[15:0],io__wdata[15:0],io__wdata[15:0],io__wdata[15:0]}; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 311:22]
  wire [63:0] _reqWdata_T_8 = {io__wdata[31:0],io__wdata[31:0]}; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 312:22]
  wire  _reqWdata_T_9 = 2'h0 == io__in_bits_func[1:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _reqWdata_T_10 = 2'h1 == io__in_bits_func[1:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _reqWdata_T_11 = 2'h2 == io__in_bits_func[1:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _reqWdata_T_12 = 2'h3 == io__in_bits_func[1:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _reqWdata_T_13 = _reqWdata_T_9 ? _reqWdata_T_3 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _reqWdata_T_14 = _reqWdata_T_10 ? _reqWdata_T_6 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _reqWdata_T_15 = _reqWdata_T_11 ? _reqWdata_T_8 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _reqWdata_T_16 = _reqWdata_T_12 ? io__wdata : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _reqWdata_T_17 = _reqWdata_T_13 | _reqWdata_T_14; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _reqWdata_T_18 = _reqWdata_T_17 | _reqWdata_T_15; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _reqWmask_T_5 = _reqWdata_T_10 ? 2'h3 : 2'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _reqWmask_T_6 = _reqWdata_T_11 ? 4'hf : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] _reqWmask_T_7 = _reqWdata_T_12 ? 8'hff : 8'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _GEN_13 = {{1'd0}, _reqWdata_T_9}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _reqWmask_T_8 = _GEN_13 | _reqWmask_T_5; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _GEN_14 = {{2'd0}, _reqWmask_T_8}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _reqWmask_T_9 = _GEN_14 | _reqWmask_T_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] _GEN_15 = {{4'd0}, _reqWmask_T_9}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] _reqWmask_T_10 = _GEN_15 | _reqWmask_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [14:0] _GEN_0 = {{7'd0}, _reqWmask_T_10}; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 306:8]
  wire [14:0] reqWmask = _GEN_0 << io__in_bits_src1[2:0]; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 306:8]
  wire  _io_out_valid_T_8 = partialLoad ? state == 2'h3 : _T_16 & state == 2'h2; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 382:114]
  reg [63:0] rdataLatch; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 388:27]
  wire  _rdataSel64_T_9 = 3'h0 == addrLatch[2:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataSel64_T_10 = 3'h1 == addrLatch[2:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataSel64_T_11 = 3'h2 == addrLatch[2:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataSel64_T_12 = 3'h3 == addrLatch[2:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataSel64_T_13 = 3'h4 == addrLatch[2:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataSel64_T_14 = 3'h5 == addrLatch[2:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataSel64_T_15 = 3'h6 == addrLatch[2:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataSel64_T_16 = 3'h7 == addrLatch[2:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdataSel64_T_17 = _rdataSel64_T_9 ? rdataLatch : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [55:0] _rdataSel64_T_18 = _rdataSel64_T_10 ? rdataLatch[63:8] : 56'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [47:0] _rdataSel64_T_19 = _rdataSel64_T_11 ? rdataLatch[63:16] : 48'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [39:0] _rdataSel64_T_20 = _rdataSel64_T_12 ? rdataLatch[63:24] : 40'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdataSel64_T_21 = _rdataSel64_T_13 ? rdataLatch[63:32] : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [23:0] _rdataSel64_T_22 = _rdataSel64_T_14 ? rdataLatch[63:40] : 24'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [15:0] _rdataSel64_T_23 = _rdataSel64_T_15 ? rdataLatch[63:48] : 16'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] _rdataSel64_T_24 = _rdataSel64_T_16 ? rdataLatch[63:56] : 8'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_16 = {{8'd0}, _rdataSel64_T_18}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataSel64_T_25 = _rdataSel64_T_17 | _GEN_16; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_17 = {{16'd0}, _rdataSel64_T_19}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataSel64_T_26 = _rdataSel64_T_25 | _GEN_17; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_18 = {{24'd0}, _rdataSel64_T_20}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataSel64_T_27 = _rdataSel64_T_26 | _GEN_18; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_19 = {{32'd0}, _rdataSel64_T_21}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataSel64_T_28 = _rdataSel64_T_27 | _GEN_19; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_20 = {{40'd0}, _rdataSel64_T_22}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataSel64_T_29 = _rdataSel64_T_28 | _GEN_20; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_21 = {{48'd0}, _rdataSel64_T_23}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataSel64_T_30 = _rdataSel64_T_29 | _GEN_21; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_22 = {{56'd0}, _rdataSel64_T_24}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] rdataSel64 = _rdataSel64_T_30 | _GEN_22; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  rdataPartialLoad_signBit = rdataSel64[7]; // @[src/main/scala/utils/BitUtils.scala 39:20]
  wire [55:0] _rdataPartialLoad_T_2 = rdataPartialLoad_signBit ? 56'hffffffffffffff : 56'h0; // @[src/main/scala/utils/BitUtils.scala 40:46]
  wire [63:0] _rdataPartialLoad_T_3 = {_rdataPartialLoad_T_2,rdataSel64[7:0]}; // @[src/main/scala/utils/BitUtils.scala 40:41]
  wire  rdataPartialLoad_signBit_1 = rdataSel64[15]; // @[src/main/scala/utils/BitUtils.scala 39:20]
  wire [47:0] _rdataPartialLoad_T_6 = rdataPartialLoad_signBit_1 ? 48'hffffffffffff : 48'h0; // @[src/main/scala/utils/BitUtils.scala 40:46]
  wire [63:0] _rdataPartialLoad_T_7 = {_rdataPartialLoad_T_6,rdataSel64[15:0]}; // @[src/main/scala/utils/BitUtils.scala 40:41]
  wire  rdataPartialLoad_signBit_2 = rdataSel64[31]; // @[src/main/scala/utils/BitUtils.scala 39:20]
  wire [31:0] _rdataPartialLoad_T_10 = rdataPartialLoad_signBit_2 ? 32'hffffffff : 32'h0; // @[src/main/scala/utils/BitUtils.scala 40:46]
  wire [63:0] _rdataPartialLoad_T_11 = {_rdataPartialLoad_T_10,rdataSel64[31:0]}; // @[src/main/scala/utils/BitUtils.scala 40:41]
  wire [63:0] _rdataPartialLoad_T_13 = {56'h0,rdataSel64[7:0]}; // @[src/main/scala/utils/BitUtils.scala 47:41]
  wire [63:0] _rdataPartialLoad_T_15 = {48'h0,rdataSel64[15:0]}; // @[src/main/scala/utils/BitUtils.scala 47:41]
  wire [63:0] _rdataPartialLoad_T_17 = {32'h0,rdataSel64[31:0]}; // @[src/main/scala/utils/BitUtils.scala 47:41]
  wire  _rdataPartialLoad_T_18 = 7'h0 == io__in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataPartialLoad_T_19 = 7'h1 == io__in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataPartialLoad_T_20 = 7'h2 == io__in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataPartialLoad_T_21 = 7'h4 == io__in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataPartialLoad_T_22 = 7'h5 == io__in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataPartialLoad_T_23 = 7'h6 == io__in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdataPartialLoad_T_24 = _rdataPartialLoad_T_18 ? _rdataPartialLoad_T_3 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_25 = _rdataPartialLoad_T_19 ? _rdataPartialLoad_T_7 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_26 = _rdataPartialLoad_T_20 ? _rdataPartialLoad_T_11 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_27 = _rdataPartialLoad_T_21 ? _rdataPartialLoad_T_13 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_28 = _rdataPartialLoad_T_22 ? _rdataPartialLoad_T_15 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_29 = _rdataPartialLoad_T_23 ? _rdataPartialLoad_T_17 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_30 = _rdataPartialLoad_T_24 | _rdataPartialLoad_T_25; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_31 = _rdataPartialLoad_T_30 | _rdataPartialLoad_T_26; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_32 = _rdataPartialLoad_T_31 | _rdataPartialLoad_T_27; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_33 = _rdataPartialLoad_T_32 | _rdataPartialLoad_T_28; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] rdataPartialLoad = _rdataPartialLoad_T_33 | _rdataPartialLoad_T_29; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _addrAligned_T_2 = ~io__in_bits_src1[0]; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 416:27]
  wire  _addrAligned_T_4 = io__in_bits_src1[1:0] == 2'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 417:29]
  wire  _addrAligned_T_6 = io__in_bits_src1[2:0] == 3'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 418:29]
  wire  addrAligned = _reqWdata_T_9 | _reqWdata_T_10 & _addrAligned_T_2 | _reqWdata_T_11 & _addrAligned_T_4 |
    _reqWdata_T_12 & _addrAligned_T_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_loadAddrMisaligned_T_4 = ~addrAligned; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 429:60]
  wire  _T_58 = ~io__dmem_req_bits_cmd[0] & ~io__dmem_req_bits_cmd[3]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:26]
  wire  _T_59 = io__dmem_req_valid & _T_58; // @[src/main/scala/bus/simplebus/SimpleBus.scala 104:29]
  wire  _T_61 = _T_59 & _T_6; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 438:39]
  reg  r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_9 = _T_59 | r; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  _T_70 = io__dmem_req_valid & io__dmem_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 103:29]
  reg  r_1; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_11 = _T_70 | r_1; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  assign io__out_valid = io__loadAddrMisaligned | io__storeAddrMisaligned | _io_out_valid_T_8; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 382:22]
  assign io__out_bits = partialLoad ? rdataPartialLoad : io__dmem_resp_bits_rdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 421:21]
  assign io__dmem_req_valid = io__in_valid & state == 2'h0 & ~io__loadAddrMisaligned & ~io__storeAddrMisaligned; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 379:75]
  assign io__dmem_req_bits_addr = io__in_bits_src1[38:0]; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 370:68]
  assign io__dmem_req_bits_size = {{1'd0}, io__in_bits_func[1:0]}; // @[src/main/scala/bus/simplebus/SimpleBus.scala 66:15]
  assign io__dmem_req_bits_cmd = {{3'd0}, isStore}; // @[src/main/scala/bus/simplebus/SimpleBus.scala 65:14]
  assign io__dmem_req_bits_wmask = reqWmask[7:0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 68:16]
  assign io__dmem_req_bits_wdata = _reqWdata_T_18 | _reqWdata_T_16; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io__dmem_resp_ready = 1'h1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 380:19]
  assign io__isMMIO = 1'h0;
  assign io__loadAddrMisaligned = io__in_valid & _partialLoad_T & ~ISAMO2 & ~addrAligned; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 429:57]
  assign io__storeAddrMisaligned = io__in_valid & (isStore | ISAMO2) & _io_loadAddrMisaligned_T_4; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 430:57]
  assign io_in_bits_src1 = io__in_bits_src1;
  always @(posedge clock) begin
    addrLatch <= io__in_bits_src1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 333:26]
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 338:22]
      state <= 2'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 338:22]
    end else if (2'h0 == state) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 351:18]
      if (_T_6) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 354:43]
        state <= 2'h2; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 354:51]
      end
    end else if (!(2'h1 == state)) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 351:18]
      if (2'h2 == state) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 351:18]
        state <= _GEN_4;
      end else begin
        state <= _GEN_5;
      end
    end
    rdataLatch <= io__dmem_resp_bits_rdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 388:27]
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (_T_16) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      r <= _GEN_9;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r_1 <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (_T_16) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      r_1 <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      r_1 <= _GEN_11;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io__in_bits_src1[63:38] == 26'h0)) begin
          $fwrite(32'h80000002,
            "Assumption failed\n    at UnpipelinedLSU.scala:331 assume(addr(XLEN - 1, VAddrBits - 1) === 0.U)\n"); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 331:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  addrLatch = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[1:0];
  _RAND_2 = {2{`RANDOM}};
  rdataLatch = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  r = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  r_1 = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assume(io__in_bits_src1[63:38] == 26'h0); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 331:9]
    end
  end
endmodule
module AtomALU(
  input  [63:0] io_src1, // @[src/main/scala/nutcore/backend/fu/LSU.scala 171:14]
  input  [63:0] io_src2, // @[src/main/scala/nutcore/backend/fu/LSU.scala 171:14]
  input  [6:0]  io_func, // @[src/main/scala/nutcore/backend/fu/LSU.scala 171:14]
  input         io_isWordOp, // @[src/main/scala/nutcore/backend/fu/LSU.scala 171:14]
  output [63:0] io_result // @[src/main/scala/nutcore/backend/fu/LSU.scala 171:14]
);
  wire  isAdderSub = ~io_func[6]; // @[src/main/scala/nutcore/backend/fu/LSU.scala 184:20]
  wire [63:0] _adderRes_T_1 = isAdderSub ? 64'hffffffffffffffff : 64'h0; // @[src/main/scala/nutcore/backend/fu/LSU.scala 185:39]
  wire [63:0] _adderRes_T_2 = io_src2 ^ _adderRes_T_1; // @[src/main/scala/nutcore/backend/fu/LSU.scala 185:33]
  wire [64:0] _adderRes_T_3 = io_src1 + _adderRes_T_2; // @[src/main/scala/nutcore/backend/fu/LSU.scala 185:24]
  wire [64:0] _GEN_0 = {{64'd0}, isAdderSub}; // @[src/main/scala/nutcore/backend/fu/LSU.scala 185:60]
  wire [64:0] adderRes = _adderRes_T_3 + _GEN_0; // @[src/main/scala/nutcore/backend/fu/LSU.scala 185:60]
  wire [63:0] xorRes = io_src1 ^ io_src2; // @[src/main/scala/nutcore/backend/fu/LSU.scala 186:21]
  wire  sltu = ~adderRes[64]; // @[src/main/scala/nutcore/backend/fu/LSU.scala 187:14]
  wire  slt = xorRes[63] ^ sltu; // @[src/main/scala/nutcore/backend/fu/LSU.scala 188:28]
  wire [63:0] _res_T_1 = io_src1 & io_src2; // @[src/main/scala/nutcore/backend/fu/LSU.scala 194:32]
  wire [63:0] _res_T_2 = io_src1 | io_src2; // @[src/main/scala/nutcore/backend/fu/LSU.scala 195:32]
  wire [63:0] _res_T_4 = slt ? io_src1 : io_src2; // @[src/main/scala/nutcore/backend/fu/LSU.scala 196:29]
  wire [63:0] _res_T_6 = slt ? io_src2 : io_src1; // @[src/main/scala/nutcore/backend/fu/LSU.scala 197:29]
  wire [63:0] _res_T_8 = sltu ? io_src1 : io_src2; // @[src/main/scala/nutcore/backend/fu/LSU.scala 198:29]
  wire [63:0] _res_T_10 = sltu ? io_src2 : io_src1; // @[src/main/scala/nutcore/backend/fu/LSU.scala 199:29]
  wire [64:0] _res_T_12 = 6'h22 == io_func[5:0] ? {{1'd0}, io_src2} : adderRes; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_14 = 6'h24 == io_func[5:0] ? {{1'd0}, xorRes} : _res_T_12; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_16 = 6'h25 == io_func[5:0] ? {{1'd0}, _res_T_1} : _res_T_14; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_18 = 6'h26 == io_func[5:0] ? {{1'd0}, _res_T_2} : _res_T_16; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_20 = 6'h37 == io_func[5:0] ? {{1'd0}, _res_T_4} : _res_T_18; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_22 = 6'h30 == io_func[5:0] ? {{1'd0}, _res_T_6} : _res_T_20; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_24 = 6'h31 == io_func[5:0] ? {{1'd0}, _res_T_8} : _res_T_22; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] res = 6'h32 == io_func[5:0] ? {{1'd0}, _res_T_10} : _res_T_24; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  io_result_signBit = res[31]; // @[src/main/scala/utils/BitUtils.scala 39:20]
  wire [31:0] _io_result_T_2 = io_result_signBit ? 32'hffffffff : 32'h0; // @[src/main/scala/utils/BitUtils.scala 40:46]
  wire [63:0] _io_result_T_3 = {_io_result_T_2,res[31:0]}; // @[src/main/scala/utils/BitUtils.scala 40:41]
  assign io_result = io_isWordOp ? _io_result_T_3 : res[63:0]; // @[src/main/scala/nutcore/backend/fu/LSU.scala 202:20]
endmodule
module UnpipelinedLSU(
  input         clock,
  input         reset,
  input         io__in_valid, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 37:14]
  input  [63:0] io__in_bits_src1, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 37:14]
  input  [63:0] io__in_bits_src2, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 37:14]
  input  [6:0]  io__in_bits_func, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 37:14]
  input         io__out_ready, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 37:14]
  output        io__out_valid, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 37:14]
  output [63:0] io__out_bits, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 37:14]
  input  [63:0] io__wdata, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 37:14]
  input  [31:0] io__instr, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 37:14]
  input         io__dmem_req_ready, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 37:14]
  output        io__dmem_req_valid, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 37:14]
  output [38:0] io__dmem_req_bits_addr, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 37:14]
  output [2:0]  io__dmem_req_bits_size, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 37:14]
  output [3:0]  io__dmem_req_bits_cmd, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 37:14]
  output [7:0]  io__dmem_req_bits_wmask, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 37:14]
  output [63:0] io__dmem_req_bits_wdata, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 37:14]
  input         io__dmem_resp_valid, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 37:14]
  input  [63:0] io__dmem_resp_bits_rdata, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 37:14]
  output        io__loadAddrMisaligned, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 37:14]
  output        io__storeAddrMisaligned, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 37:14]
  output        setLr_0,
  output [63:0] io_in_bits_src1,
  output [63:0] setLrAddr_0,
  output        setLrVal_0,
  input  [63:0] lr_addr
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  lsExecUnit_clock; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_reset; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__in_valid; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire [63:0] lsExecUnit_io__in_bits_src1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire [6:0] lsExecUnit_io__in_bits_func; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__out_ready; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__out_valid; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire [63:0] lsExecUnit_io__out_bits; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire [63:0] lsExecUnit_io__wdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__dmem_req_ready; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__dmem_req_valid; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire [38:0] lsExecUnit_io__dmem_req_bits_addr; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire [2:0] lsExecUnit_io__dmem_req_bits_size; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire [3:0] lsExecUnit_io__dmem_req_bits_cmd; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire [7:0] lsExecUnit_io__dmem_req_bits_wmask; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire [63:0] lsExecUnit_io__dmem_req_bits_wdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__dmem_resp_ready; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__dmem_resp_valid; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire [63:0] lsExecUnit_io__dmem_resp_bits_rdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__isMMIO; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__loadAddrMisaligned; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__storeAddrMisaligned; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_ISAMO2; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire [63:0] lsExecUnit_io_in_bits_src1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
  wire [63:0] atomALU_io_src1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 98:25]
  wire [63:0] atomALU_io_src2; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 98:25]
  wire [6:0] atomALU_io_func; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 98:25]
  wire  atomALU_io_isWordOp; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 98:25]
  wire [63:0] atomALU_io_result; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 98:25]
  wire  atomReq = io__in_valid & io__in_bits_func[5]; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 53:26]
  wire  _amoReq_T_1 = io__in_bits_func == 7'h20; // @[src/main/scala/nutcore/backend/fu/LSU.scala 57:37]
  wire  _amoReq_T_4 = io__in_bits_func == 7'h21; // @[src/main/scala/nutcore/backend/fu/LSU.scala 58:37]
  wire  _amoReq_T_6 = io__in_bits_func[5] & ~_amoReq_T_1 & ~_amoReq_T_4; // @[src/main/scala/nutcore/backend/fu/LSU.scala 59:61]
  wire  amoReq = io__in_valid & _amoReq_T_6; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 54:26]
  wire  lrReq = io__in_valid & _amoReq_T_1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 55:25]
  wire  scReq = io__in_valid & _amoReq_T_4; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 56:25]
  wire [2:0] funct3 = io__instr[14:12]; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 64:26]
  wire  scInvalid = ~(io__in_bits_src1 == lr_addr) & scReq; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 81:40]
  reg [2:0] state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 95:24]
  reg [63:0] atomMemReg; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 96:25]
  reg [63:0] atomRegReg; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 97:25]
  wire  _T = 3'h0 == state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20]
  wire  _lsExecUnit_io_in_valid_T = ~atomReq; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 141:56]
  wire [63:0] _lsExecUnit_io_in_bits_src1_T_1 = io__in_bits_src1 + io__in_bits_src2; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 143:46]
  wire  _io_in_ready_T_1 = lsExecUnit_io__out_ready & lsExecUnit_io__out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [2:0] _GEN_1 = amoReq ? 3'h5 : 3'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 149:17 152:{21,28}]
  wire [2:0] _GEN_2 = lrReq ? 3'h3 : _GEN_1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 153:{20,27}]
  wire [2:0] _state_T = scInvalid ? 3'h0 : 3'h4; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 154:33]
  wire  _T_1 = 3'h1 == state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20]
  wire [2:0] _GEN_4 = io__out_valid ? 3'h0 : state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 168:{26,33} 95:24]
  wire [1:0] _lsExecUnit_io_in_bits_func_T = funct3[0] ? 2'h3 : 2'h2; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 188:42]
  wire [2:0] _GEN_5 = _io_in_ready_T_1 ? 3'h6 : state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 192:37 193:17 95:24]
  wire [3:0] _lsExecUnit_io_in_bits_func_T_1 = funct3[0] ? 4'hb : 4'ha; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 219:42]
  wire [2:0] _GEN_6 = _io_in_ready_T_1 ? 3'h0 : state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 223:37 224:17 95:24]
  wire [63:0] _GEN_11 = io__in_bits_src1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 245:36]
  wire  _GEN_14 = 3'h4 == state & _io_in_ready_T_1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 126:32 249:36]
  wire [2:0] _GEN_16 = 3'h4 == state ? _GEN_6 : state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 95:24]
  wire  _GEN_17 = 3'h3 == state | 3'h4 == state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 229:36]
  wire [3:0] _GEN_20 = 3'h3 == state ? {{2'd0}, _lsExecUnit_io_in_bits_func_T} : _lsExecUnit_io_in_bits_func_T_1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 233:36]
  wire  _GEN_22 = 3'h3 == state ? _io_in_ready_T_1 : _GEN_14; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 235:36]
  wire [2:0] _GEN_24 = 3'h3 == state ? _GEN_6 : _GEN_16; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20]
  wire  _GEN_25 = 3'h7 == state | _GEN_17; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 215:36]
  wire [3:0] _GEN_28 = 3'h7 == state ? _lsExecUnit_io_in_bits_func_T_1 : _GEN_20; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 219:36]
  wire [63:0] _GEN_29 = 3'h7 == state ? atomMemReg : io__wdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 220:36]
  wire  _GEN_30 = 3'h7 == state ? _io_in_ready_T_1 : _GEN_22; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 221:36]
  wire [2:0] _GEN_32 = 3'h7 == state ? _GEN_6 : _GEN_24; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20]
  wire  _GEN_33 = 3'h6 == state ? 1'h0 : _GEN_25; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 201:36]
  wire  _GEN_34 = 3'h6 == state ? 1'h0 : 1'h1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 202:36]
  wire  _GEN_38 = 3'h6 == state ? 1'h0 : _GEN_30; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 207:36]
  wire [2:0] _GEN_40 = 3'h6 == state ? 3'h7 : _GEN_32; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 209:15]
  wire  _GEN_42 = 3'h5 == state | _GEN_33; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 184:36]
  wire  _GEN_43 = 3'h5 == state | _GEN_34; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 185:36]
  wire [3:0] _GEN_45 = 3'h5 == state ? {{2'd0}, _lsExecUnit_io_in_bits_func_T} : _GEN_28; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 188:36]
  wire  _GEN_47 = 3'h5 == state ? 1'h0 : _GEN_38; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 190:36]
  wire [2:0] _GEN_49 = 3'h5 == state ? _GEN_5 : _GEN_40; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20]
  wire  _GEN_52 = 3'h1 == state | _GEN_42; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 159:36]
  wire  _GEN_53 = 3'h1 == state | _GEN_43; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 160:36]
  wire [6:0] _GEN_55 = 3'h1 == state ? io__in_bits_func : {{3'd0}, _GEN_45}; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 163:36]
  wire [63:0] _GEN_56 = 3'h1 == state ? io__wdata : _GEN_29; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 164:36]
  wire  _GEN_58 = 3'h1 == state ? lsExecUnit_io__out_valid : _GEN_47; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 166:36]
  wire  _GEN_68 = 3'h0 == state ? lsExecUnit_io__out_valid | scInvalid : _GEN_58; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 148:38]
  wire [63:0] _io_out_bits_T_1 = state == 3'h7 ? atomRegReg : lsExecUnit_io__out_bits; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 275:45]
  wire  setLr = io__out_valid & (lrReq | scReq); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 270:26]
  wire  setLrVal = lrReq; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 55:25]
  wire [63:0] setLrAddr = io__in_bits_src1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 272:15 72:25]
  LSExecUnit lsExecUnit ( // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 47:28]
    .clock(lsExecUnit_clock),
    .reset(lsExecUnit_reset),
    .io__in_valid(lsExecUnit_io__in_valid),
    .io__in_bits_src1(lsExecUnit_io__in_bits_src1),
    .io__in_bits_func(lsExecUnit_io__in_bits_func),
    .io__out_ready(lsExecUnit_io__out_ready),
    .io__out_valid(lsExecUnit_io__out_valid),
    .io__out_bits(lsExecUnit_io__out_bits),
    .io__wdata(lsExecUnit_io__wdata),
    .io__dmem_req_ready(lsExecUnit_io__dmem_req_ready),
    .io__dmem_req_valid(lsExecUnit_io__dmem_req_valid),
    .io__dmem_req_bits_addr(lsExecUnit_io__dmem_req_bits_addr),
    .io__dmem_req_bits_size(lsExecUnit_io__dmem_req_bits_size),
    .io__dmem_req_bits_cmd(lsExecUnit_io__dmem_req_bits_cmd),
    .io__dmem_req_bits_wmask(lsExecUnit_io__dmem_req_bits_wmask),
    .io__dmem_req_bits_wdata(lsExecUnit_io__dmem_req_bits_wdata),
    .io__dmem_resp_ready(lsExecUnit_io__dmem_resp_ready),
    .io__dmem_resp_valid(lsExecUnit_io__dmem_resp_valid),
    .io__dmem_resp_bits_rdata(lsExecUnit_io__dmem_resp_bits_rdata),
    .io__isMMIO(lsExecUnit_io__isMMIO),
    .io__loadAddrMisaligned(lsExecUnit_io__loadAddrMisaligned),
    .io__storeAddrMisaligned(lsExecUnit_io__storeAddrMisaligned),
    .ISAMO2(lsExecUnit_ISAMO2),
    .io_in_bits_src1(lsExecUnit_io_in_bits_src1)
  );
  AtomALU atomALU ( // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 98:25]
    .io_src1(atomALU_io_src1),
    .io_src2(atomALU_io_src2),
    .io_func(atomALU_io_func),
    .io_isWordOp(atomALU_io_isWordOp),
    .io_result(atomALU_io_result)
  );
  assign io__out_valid = io__loadAddrMisaligned | io__storeAddrMisaligned | _GEN_68; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 257:68 259:20]
  assign io__out_bits = scReq ? {{63'd0}, scInvalid} : _io_out_bits_T_1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 275:23]
  assign io__dmem_req_valid = lsExecUnit_io__dmem_req_valid; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 274:13]
  assign io__dmem_req_bits_addr = lsExecUnit_io__dmem_req_bits_addr; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 274:13]
  assign io__dmem_req_bits_size = lsExecUnit_io__dmem_req_bits_size; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 274:13]
  assign io__dmem_req_bits_cmd = lsExecUnit_io__dmem_req_bits_cmd; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 274:13]
  assign io__dmem_req_bits_wmask = lsExecUnit_io__dmem_req_bits_wmask; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 274:13]
  assign io__dmem_req_bits_wdata = lsExecUnit_io__dmem_req_bits_wdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 274:13]
  assign io__loadAddrMisaligned = lsExecUnit_io__loadAddrMisaligned; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 285:27]
  assign io__storeAddrMisaligned = lsExecUnit_io__storeAddrMisaligned; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 286:28]
  assign setLr_0 = setLr;
  assign io_in_bits_src1 = lsExecUnit_io_in_bits_src1;
  assign setLrAddr_0 = _GEN_11;
  assign setLrVal_0 = setLrVal;
  assign lsExecUnit_clock = clock;
  assign lsExecUnit_reset = reset;
  assign lsExecUnit_io__in_valid = 3'h0 == state ? io__in_valid & ~atomReq : _GEN_52; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 141:38]
  assign lsExecUnit_io__in_bits_src1 = 3'h0 == state ? _lsExecUnit_io_in_bits_src1_T_1 : io__in_bits_src1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 143:38]
  assign lsExecUnit_io__in_bits_func = 3'h0 == state ? io__in_bits_func : _GEN_55; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 145:38]
  assign lsExecUnit_io__out_ready = 3'h0 == state | _GEN_53; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 142:38]
  assign lsExecUnit_io__wdata = 3'h0 == state ? io__wdata : _GEN_56; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20 146:38]
  assign lsExecUnit_io__dmem_req_ready = io__dmem_req_ready; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 274:13]
  assign lsExecUnit_io__dmem_resp_valid = io__dmem_resp_valid; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 274:13]
  assign lsExecUnit_io__dmem_resp_bits_rdata = io__dmem_resp_bits_rdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 274:13]
  assign lsExecUnit_ISAMO2 = amoReq;
  assign atomALU_io_src1 = atomMemReg; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 99:21]
  assign atomALU_io_src2 = io__wdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 100:21]
  assign atomALU_io_func = io__in_bits_func; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 101:21]
  assign atomALU_io_isWordOp = ~funct3[0]; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 66:22]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 95:24]
      state <= 3'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 95:24]
    end else if (io__loadAddrMisaligned | io__storeAddrMisaligned) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 257:68]
      state <= 3'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 258:13]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20]
      if (scReq) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 154:20]
        state <= _state_T; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 154:27]
      end else begin
        state <= _GEN_2;
      end
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20]
      state <= _GEN_4;
    end else begin
      state <= _GEN_49;
    end
    if (!(3'h0 == state)) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20]
      if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20]
        if (3'h5 == state) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20]
          atomMemReg <= lsExecUnit_io__out_bits; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 196:20]
        end else if (3'h6 == state) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20]
          atomMemReg <= atomALU_io_result; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 210:20]
        end
      end
    end
    if (!(3'h0 == state)) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20]
      if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20]
        if (3'h5 == state) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 128:20]
          atomRegReg <= lsExecUnit_io__out_bits; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 197:20]
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T & _T_1 & ~reset & ~(_lsExecUnit_io_in_valid_T | ~amoReq | ~lrReq | ~scReq)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at UnpipelinedLSU.scala:167 assert(!atomReq || !amoReq || !lrReq || !scReq)\n"); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 167:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {2{`RANDOM}};
  atomMemReg = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  atomRegReg = _RAND_2[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~_T & _T_1 & ~reset) begin
      assert(_lsExecUnit_io_in_valid_T | ~amoReq | ~lrReq | ~scReq); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 167:15]
    end
  end
endmodule
module Multiplier(
  input          clock,
  input          reset,
  output         io_in_ready, // @[src/main/scala/nutcore/backend/fu/MDU.scala 53:14]
  input          io_in_valid, // @[src/main/scala/nutcore/backend/fu/MDU.scala 53:14]
  input  [64:0]  io_in_bits_0, // @[src/main/scala/nutcore/backend/fu/MDU.scala 53:14]
  input  [64:0]  io_in_bits_1, // @[src/main/scala/nutcore/backend/fu/MDU.scala 53:14]
  input          io_out_ready, // @[src/main/scala/nutcore/backend/fu/MDU.scala 53:14]
  output         io_out_valid, // @[src/main/scala/nutcore/backend/fu/MDU.scala 53:14]
  output [129:0] io_out_bits // @[src/main/scala/nutcore/backend/fu/MDU.scala 53:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [95:0] _RAND_0;
  reg [95:0] _RAND_1;
  reg [159:0] _RAND_2;
  reg [159:0] _RAND_3;
  reg [159:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  reg [64:0] mulRes_REG; // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
  reg [64:0] mulRes_REG_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
  reg [129:0] io_out_bits_REG; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
  reg [129:0] io_out_bits_REG_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
  reg [129:0] io_out_bits_REG_2; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
  reg  io_out_valid_REG; // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
  reg  io_out_valid_REG_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
  reg  io_out_valid_REG_2; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
  reg  io_out_valid_REG_3; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
  reg  busy; // @[src/main/scala/nutcore/backend/fu/MDU.scala 62:21]
  wire  _GEN_0 = io_in_valid & ~busy | busy; // @[src/main/scala/nutcore/backend/fu/MDU.scala 62:21 63:{31,38}]
  assign io_in_ready = ~busy; // @[src/main/scala/nutcore/backend/fu/MDU.scala 65:49]
  assign io_out_valid = io_out_valid_REG_3; // @[src/main/scala/nutcore/backend/fu/MDU.scala 60:16]
  assign io_out_bits = io_out_bits_REG_2; // @[src/main/scala/nutcore/backend/fu/MDU.scala 59:37]
  always @(posedge clock) begin
    mulRes_REG <= io_in_bits_0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    mulRes_REG_1 <= io_in_bits_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    io_out_bits_REG <= $signed(mulRes_REG) * $signed(mulRes_REG_1); // @[src/main/scala/nutcore/backend/fu/MDU.scala 58:49]
    io_out_bits_REG_1 <= io_out_bits_REG; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    io_out_bits_REG_2 <= io_out_bits_REG_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    io_out_valid_REG <= io_in_ready & io_in_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
    io_out_valid_REG_1 <= io_out_valid_REG; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    io_out_valid_REG_2 <= io_out_valid_REG_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    io_out_valid_REG_3 <= io_out_valid_REG_2; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 62:21]
      busy <= 1'h0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 62:21]
    end else if (io_out_valid) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 64:23]
      busy <= 1'h0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 64:30]
    end else begin
      busy <= _GEN_0;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {3{`RANDOM}};
  mulRes_REG = _RAND_0[64:0];
  _RAND_1 = {3{`RANDOM}};
  mulRes_REG_1 = _RAND_1[64:0];
  _RAND_2 = {5{`RANDOM}};
  io_out_bits_REG = _RAND_2[129:0];
  _RAND_3 = {5{`RANDOM}};
  io_out_bits_REG_1 = _RAND_3[129:0];
  _RAND_4 = {5{`RANDOM}};
  io_out_bits_REG_2 = _RAND_4[129:0];
  _RAND_5 = {1{`RANDOM}};
  io_out_valid_REG = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  io_out_valid_REG_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  io_out_valid_REG_2 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  io_out_valid_REG_3 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  busy = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Divider(
  input          clock,
  input          reset,
  output         io_in_ready, // @[src/main/scala/nutcore/backend/fu/MDU.scala 69:14]
  input          io_in_valid, // @[src/main/scala/nutcore/backend/fu/MDU.scala 69:14]
  input  [63:0]  io_in_bits_0, // @[src/main/scala/nutcore/backend/fu/MDU.scala 69:14]
  input  [63:0]  io_in_bits_1, // @[src/main/scala/nutcore/backend/fu/MDU.scala 69:14]
  input          io_sign, // @[src/main/scala/nutcore/backend/fu/MDU.scala 69:14]
  output         io_out_valid, // @[src/main/scala/nutcore/backend/fu/MDU.scala 69:14]
  output [127:0] io_out_bits // @[src/main/scala/nutcore/backend/fu/MDU.scala 69:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [159:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [95:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[src/main/scala/nutcore/backend/fu/MDU.scala 77:22]
  wire  _newReq_T_1 = io_in_ready & io_in_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  newReq = state == 3'h0 & _newReq_T_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 78:35]
  wire  divBy0 = io_in_bits_1 == 64'h0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 81:18]
  reg [128:0] shiftReg; // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
  wire [64:0] hi = shiftReg[128:64]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 84:20]
  wire [63:0] lo = shiftReg[63:0]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 85:20]
  wire  aSign = io_in_bits_0[63] & io_sign; // @[src/main/scala/nutcore/backend/fu/MDU.scala 72:24]
  wire [63:0] _T_1 = 64'h0 - io_in_bits_0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 73:16]
  wire [63:0] aVal = aSign ? _T_1 : io_in_bits_0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 73:12]
  wire  bSign = io_in_bits_1[63] & io_sign; // @[src/main/scala/nutcore/backend/fu/MDU.scala 72:24]
  wire [63:0] _T_3 = 64'h0 - io_in_bits_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 73:16]
  reg  aSignReg; // @[src/main/scala/nutcore/backend/fu/MDU.scala 89:27]
  reg  qSignReg; // @[src/main/scala/nutcore/backend/fu/MDU.scala 90:27]
  reg [63:0] bReg; // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
  wire [64:0] _aValx2Reg_T = {aVal,1'h0}; // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:32]
  reg [64:0] aValx2Reg; // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
  reg [5:0] cnt_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [31:0] canSkipShift_hi = bReg[63:32]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [31:0] canSkipShift_lo = bReg[31:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi = |canSkipShift_hi; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [15:0] canSkipShift_hi_1 = canSkipShift_hi[31:16]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [15:0] canSkipShift_lo_1 = canSkipShift_hi[15:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_1 = |canSkipShift_hi_1; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [7:0] canSkipShift_hi_2 = canSkipShift_hi_1[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] canSkipShift_lo_2 = canSkipShift_hi_1[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_2 = |canSkipShift_hi_2; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] canSkipShift_hi_3 = canSkipShift_hi_2[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_3 = canSkipShift_hi_2[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_3 = |canSkipShift_hi_3; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_3 = canSkipShift_hi_3[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_3[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_4 = canSkipShift_hi_3[3] ? 2'h3 : _canSkipShift_T_3; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_8 = canSkipShift_lo_3[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_3[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_9 = canSkipShift_lo_3[3] ? 2'h3 : _canSkipShift_T_8; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_10 = canSkipShift_useHi_3 ? _canSkipShift_T_4 : _canSkipShift_T_9; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_11 = {canSkipShift_useHi_3,_canSkipShift_T_10}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] canSkipShift_hi_4 = canSkipShift_lo_2[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_4 = canSkipShift_lo_2[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_4 = |canSkipShift_hi_4; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_15 = canSkipShift_hi_4[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_4[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_16 = canSkipShift_hi_4[3] ? 2'h3 : _canSkipShift_T_15; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_20 = canSkipShift_lo_4[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_4[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_21 = canSkipShift_lo_4[3] ? 2'h3 : _canSkipShift_T_20; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_22 = canSkipShift_useHi_4 ? _canSkipShift_T_16 : _canSkipShift_T_21; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_23 = {canSkipShift_useHi_4,_canSkipShift_T_22}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _canSkipShift_T_24 = canSkipShift_useHi_2 ? _canSkipShift_T_11 : _canSkipShift_T_23; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _canSkipShift_T_25 = {canSkipShift_useHi_2,_canSkipShift_T_24}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [7:0] canSkipShift_hi_5 = canSkipShift_lo_1[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] canSkipShift_lo_5 = canSkipShift_lo_1[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_5 = |canSkipShift_hi_5; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] canSkipShift_hi_6 = canSkipShift_hi_5[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_6 = canSkipShift_hi_5[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_6 = |canSkipShift_hi_6; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_29 = canSkipShift_hi_6[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_6[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_30 = canSkipShift_hi_6[3] ? 2'h3 : _canSkipShift_T_29; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_34 = canSkipShift_lo_6[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_6[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_35 = canSkipShift_lo_6[3] ? 2'h3 : _canSkipShift_T_34; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_36 = canSkipShift_useHi_6 ? _canSkipShift_T_30 : _canSkipShift_T_35; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_37 = {canSkipShift_useHi_6,_canSkipShift_T_36}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] canSkipShift_hi_7 = canSkipShift_lo_5[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_7 = canSkipShift_lo_5[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_7 = |canSkipShift_hi_7; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_41 = canSkipShift_hi_7[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_7[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_42 = canSkipShift_hi_7[3] ? 2'h3 : _canSkipShift_T_41; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_46 = canSkipShift_lo_7[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_7[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_47 = canSkipShift_lo_7[3] ? 2'h3 : _canSkipShift_T_46; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_48 = canSkipShift_useHi_7 ? _canSkipShift_T_42 : _canSkipShift_T_47; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_49 = {canSkipShift_useHi_7,_canSkipShift_T_48}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _canSkipShift_T_50 = canSkipShift_useHi_5 ? _canSkipShift_T_37 : _canSkipShift_T_49; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _canSkipShift_T_51 = {canSkipShift_useHi_5,_canSkipShift_T_50}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] _canSkipShift_T_52 = canSkipShift_useHi_1 ? _canSkipShift_T_25 : _canSkipShift_T_51; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [4:0] _canSkipShift_T_53 = {canSkipShift_useHi_1,_canSkipShift_T_52}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [15:0] canSkipShift_hi_8 = canSkipShift_lo[31:16]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [15:0] canSkipShift_lo_8 = canSkipShift_lo[15:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_8 = |canSkipShift_hi_8; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [7:0] canSkipShift_hi_9 = canSkipShift_hi_8[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] canSkipShift_lo_9 = canSkipShift_hi_8[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_9 = |canSkipShift_hi_9; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] canSkipShift_hi_10 = canSkipShift_hi_9[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_10 = canSkipShift_hi_9[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_10 = |canSkipShift_hi_10; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_57 = canSkipShift_hi_10[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_10[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_58 = canSkipShift_hi_10[3] ? 2'h3 : _canSkipShift_T_57; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_62 = canSkipShift_lo_10[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_10[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_63 = canSkipShift_lo_10[3] ? 2'h3 : _canSkipShift_T_62; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_64 = canSkipShift_useHi_10 ? _canSkipShift_T_58 : _canSkipShift_T_63; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_65 = {canSkipShift_useHi_10,_canSkipShift_T_64}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] canSkipShift_hi_11 = canSkipShift_lo_9[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_11 = canSkipShift_lo_9[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_11 = |canSkipShift_hi_11; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_69 = canSkipShift_hi_11[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_11[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_70 = canSkipShift_hi_11[3] ? 2'h3 : _canSkipShift_T_69; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_74 = canSkipShift_lo_11[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_11[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_75 = canSkipShift_lo_11[3] ? 2'h3 : _canSkipShift_T_74; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_76 = canSkipShift_useHi_11 ? _canSkipShift_T_70 : _canSkipShift_T_75; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_77 = {canSkipShift_useHi_11,_canSkipShift_T_76}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _canSkipShift_T_78 = canSkipShift_useHi_9 ? _canSkipShift_T_65 : _canSkipShift_T_77; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _canSkipShift_T_79 = {canSkipShift_useHi_9,_canSkipShift_T_78}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [7:0] canSkipShift_hi_12 = canSkipShift_lo_8[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] canSkipShift_lo_12 = canSkipShift_lo_8[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_12 = |canSkipShift_hi_12; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] canSkipShift_hi_13 = canSkipShift_hi_12[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_13 = canSkipShift_hi_12[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_13 = |canSkipShift_hi_13; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_83 = canSkipShift_hi_13[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_13[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_84 = canSkipShift_hi_13[3] ? 2'h3 : _canSkipShift_T_83; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_88 = canSkipShift_lo_13[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_13[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_89 = canSkipShift_lo_13[3] ? 2'h3 : _canSkipShift_T_88; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_90 = canSkipShift_useHi_13 ? _canSkipShift_T_84 : _canSkipShift_T_89; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_91 = {canSkipShift_useHi_13,_canSkipShift_T_90}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] canSkipShift_hi_14 = canSkipShift_lo_12[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_14 = canSkipShift_lo_12[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_14 = |canSkipShift_hi_14; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_95 = canSkipShift_hi_14[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_14[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_96 = canSkipShift_hi_14[3] ? 2'h3 : _canSkipShift_T_95; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_100 = canSkipShift_lo_14[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_14[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_101 = canSkipShift_lo_14[3] ? 2'h3 : _canSkipShift_T_100; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_102 = canSkipShift_useHi_14 ? _canSkipShift_T_96 : _canSkipShift_T_101; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_103 = {canSkipShift_useHi_14,_canSkipShift_T_102}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _canSkipShift_T_104 = canSkipShift_useHi_12 ? _canSkipShift_T_91 : _canSkipShift_T_103; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _canSkipShift_T_105 = {canSkipShift_useHi_12,_canSkipShift_T_104}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] _canSkipShift_T_106 = canSkipShift_useHi_8 ? _canSkipShift_T_79 : _canSkipShift_T_105; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [4:0] _canSkipShift_T_107 = {canSkipShift_useHi_8,_canSkipShift_T_106}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [4:0] _canSkipShift_T_108 = canSkipShift_useHi ? _canSkipShift_T_53 : _canSkipShift_T_107; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [5:0] _canSkipShift_T_109 = {canSkipShift_useHi,_canSkipShift_T_108}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [6:0] _GEN_18 = {{1'd0}, _canSkipShift_T_109}; // @[src/main/scala/nutcore/backend/fu/MDU.scala 105:31]
  wire [6:0] _canSkipShift_T_110 = 7'h40 | _GEN_18; // @[src/main/scala/nutcore/backend/fu/MDU.scala 105:31]
  wire  canSkipShift_hi_15 = aValx2Reg[64]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [63:0] canSkipShift_lo_15 = aValx2Reg[63:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_15 = |canSkipShift_hi_15; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [31:0] canSkipShift_hi_16 = canSkipShift_lo_15[63:32]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [31:0] canSkipShift_lo_16 = canSkipShift_lo_15[31:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_16 = |canSkipShift_hi_16; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [15:0] canSkipShift_hi_17 = canSkipShift_hi_16[31:16]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [15:0] canSkipShift_lo_17 = canSkipShift_hi_16[15:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_17 = |canSkipShift_hi_17; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [7:0] canSkipShift_hi_18 = canSkipShift_hi_17[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] canSkipShift_lo_18 = canSkipShift_hi_17[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_18 = |canSkipShift_hi_18; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] canSkipShift_hi_19 = canSkipShift_hi_18[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_19 = canSkipShift_hi_18[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_19 = |canSkipShift_hi_19; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_114 = canSkipShift_hi_19[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_19[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_115 = canSkipShift_hi_19[3] ? 2'h3 : _canSkipShift_T_114; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_119 = canSkipShift_lo_19[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_19[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_120 = canSkipShift_lo_19[3] ? 2'h3 : _canSkipShift_T_119; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_121 = canSkipShift_useHi_19 ? _canSkipShift_T_115 : _canSkipShift_T_120; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_122 = {canSkipShift_useHi_19,_canSkipShift_T_121}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] canSkipShift_hi_20 = canSkipShift_lo_18[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_20 = canSkipShift_lo_18[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_20 = |canSkipShift_hi_20; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_126 = canSkipShift_hi_20[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_20[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_127 = canSkipShift_hi_20[3] ? 2'h3 : _canSkipShift_T_126; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_131 = canSkipShift_lo_20[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_20[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_132 = canSkipShift_lo_20[3] ? 2'h3 : _canSkipShift_T_131; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_133 = canSkipShift_useHi_20 ? _canSkipShift_T_127 : _canSkipShift_T_132; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_134 = {canSkipShift_useHi_20,_canSkipShift_T_133}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _canSkipShift_T_135 = canSkipShift_useHi_18 ? _canSkipShift_T_122 : _canSkipShift_T_134; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _canSkipShift_T_136 = {canSkipShift_useHi_18,_canSkipShift_T_135}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [7:0] canSkipShift_hi_21 = canSkipShift_lo_17[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] canSkipShift_lo_21 = canSkipShift_lo_17[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_21 = |canSkipShift_hi_21; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] canSkipShift_hi_22 = canSkipShift_hi_21[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_22 = canSkipShift_hi_21[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_22 = |canSkipShift_hi_22; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_140 = canSkipShift_hi_22[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_22[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_141 = canSkipShift_hi_22[3] ? 2'h3 : _canSkipShift_T_140; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_145 = canSkipShift_lo_22[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_22[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_146 = canSkipShift_lo_22[3] ? 2'h3 : _canSkipShift_T_145; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_147 = canSkipShift_useHi_22 ? _canSkipShift_T_141 : _canSkipShift_T_146; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_148 = {canSkipShift_useHi_22,_canSkipShift_T_147}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] canSkipShift_hi_23 = canSkipShift_lo_21[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_23 = canSkipShift_lo_21[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_23 = |canSkipShift_hi_23; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_152 = canSkipShift_hi_23[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_23[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_153 = canSkipShift_hi_23[3] ? 2'h3 : _canSkipShift_T_152; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_157 = canSkipShift_lo_23[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_23[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_158 = canSkipShift_lo_23[3] ? 2'h3 : _canSkipShift_T_157; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_159 = canSkipShift_useHi_23 ? _canSkipShift_T_153 : _canSkipShift_T_158; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_160 = {canSkipShift_useHi_23,_canSkipShift_T_159}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _canSkipShift_T_161 = canSkipShift_useHi_21 ? _canSkipShift_T_148 : _canSkipShift_T_160; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _canSkipShift_T_162 = {canSkipShift_useHi_21,_canSkipShift_T_161}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] _canSkipShift_T_163 = canSkipShift_useHi_17 ? _canSkipShift_T_136 : _canSkipShift_T_162; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [4:0] _canSkipShift_T_164 = {canSkipShift_useHi_17,_canSkipShift_T_163}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [15:0] canSkipShift_hi_24 = canSkipShift_lo_16[31:16]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [15:0] canSkipShift_lo_24 = canSkipShift_lo_16[15:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_24 = |canSkipShift_hi_24; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [7:0] canSkipShift_hi_25 = canSkipShift_hi_24[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] canSkipShift_lo_25 = canSkipShift_hi_24[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_25 = |canSkipShift_hi_25; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] canSkipShift_hi_26 = canSkipShift_hi_25[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_26 = canSkipShift_hi_25[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_26 = |canSkipShift_hi_26; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_168 = canSkipShift_hi_26[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_26[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_169 = canSkipShift_hi_26[3] ? 2'h3 : _canSkipShift_T_168; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_173 = canSkipShift_lo_26[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_26[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_174 = canSkipShift_lo_26[3] ? 2'h3 : _canSkipShift_T_173; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_175 = canSkipShift_useHi_26 ? _canSkipShift_T_169 : _canSkipShift_T_174; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_176 = {canSkipShift_useHi_26,_canSkipShift_T_175}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] canSkipShift_hi_27 = canSkipShift_lo_25[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_27 = canSkipShift_lo_25[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_27 = |canSkipShift_hi_27; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_180 = canSkipShift_hi_27[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_27[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_181 = canSkipShift_hi_27[3] ? 2'h3 : _canSkipShift_T_180; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_185 = canSkipShift_lo_27[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_27[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_186 = canSkipShift_lo_27[3] ? 2'h3 : _canSkipShift_T_185; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_187 = canSkipShift_useHi_27 ? _canSkipShift_T_181 : _canSkipShift_T_186; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_188 = {canSkipShift_useHi_27,_canSkipShift_T_187}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _canSkipShift_T_189 = canSkipShift_useHi_25 ? _canSkipShift_T_176 : _canSkipShift_T_188; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _canSkipShift_T_190 = {canSkipShift_useHi_25,_canSkipShift_T_189}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [7:0] canSkipShift_hi_28 = canSkipShift_lo_24[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] canSkipShift_lo_28 = canSkipShift_lo_24[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_28 = |canSkipShift_hi_28; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] canSkipShift_hi_29 = canSkipShift_hi_28[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_29 = canSkipShift_hi_28[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_29 = |canSkipShift_hi_29; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_194 = canSkipShift_hi_29[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_29[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_195 = canSkipShift_hi_29[3] ? 2'h3 : _canSkipShift_T_194; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_199 = canSkipShift_lo_29[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_29[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_200 = canSkipShift_lo_29[3] ? 2'h3 : _canSkipShift_T_199; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_201 = canSkipShift_useHi_29 ? _canSkipShift_T_195 : _canSkipShift_T_200; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_202 = {canSkipShift_useHi_29,_canSkipShift_T_201}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] canSkipShift_hi_30 = canSkipShift_lo_28[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_30 = canSkipShift_lo_28[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_30 = |canSkipShift_hi_30; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_206 = canSkipShift_hi_30[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_30[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_207 = canSkipShift_hi_30[3] ? 2'h3 : _canSkipShift_T_206; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_211 = canSkipShift_lo_30[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_30[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_212 = canSkipShift_lo_30[3] ? 2'h3 : _canSkipShift_T_211; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_213 = canSkipShift_useHi_30 ? _canSkipShift_T_207 : _canSkipShift_T_212; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_214 = {canSkipShift_useHi_30,_canSkipShift_T_213}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _canSkipShift_T_215 = canSkipShift_useHi_28 ? _canSkipShift_T_202 : _canSkipShift_T_214; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _canSkipShift_T_216 = {canSkipShift_useHi_28,_canSkipShift_T_215}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] _canSkipShift_T_217 = canSkipShift_useHi_24 ? _canSkipShift_T_190 : _canSkipShift_T_216; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [4:0] _canSkipShift_T_218 = {canSkipShift_useHi_24,_canSkipShift_T_217}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [4:0] _canSkipShift_T_219 = canSkipShift_useHi_16 ? _canSkipShift_T_164 : _canSkipShift_T_218; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [5:0] _canSkipShift_T_220 = {canSkipShift_useHi_16,_canSkipShift_T_219}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [5:0] _canSkipShift_T_221 = canSkipShift_useHi_15 ? 6'h0 : _canSkipShift_T_220; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [6:0] _canSkipShift_T_222 = {canSkipShift_useHi_15,_canSkipShift_T_221}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [6:0] canSkipShift = _canSkipShift_T_110 - _canSkipShift_T_222; // @[src/main/scala/nutcore/backend/fu/MDU.scala 105:45]
  wire [6:0] _value_T_1 = canSkipShift >= 7'h3f ? 7'h3f : canSkipShift; // @[src/main/scala/nutcore/backend/fu/MDU.scala 109:38]
  wire [6:0] _value_T_2 = divBy0 ? 7'h0 : _value_T_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 109:21]
  wire [127:0] _GEN_0 = {{63'd0}, aValx2Reg}; // @[src/main/scala/nutcore/backend/fu/MDU.scala 112:27]
  wire [127:0] _shiftReg_T = _GEN_0 << cnt_value; // @[src/main/scala/nutcore/backend/fu/MDU.scala 112:27]
  wire [64:0] _GEN_19 = {{1'd0}, bReg}; // @[src/main/scala/nutcore/backend/fu/MDU.scala 115:28]
  wire  enough = hi >= _GEN_19; // @[src/main/scala/nutcore/backend/fu/MDU.scala 115:28]
  wire [64:0] _shiftReg_T_2 = hi - _GEN_19; // @[src/main/scala/nutcore/backend/fu/MDU.scala 116:36]
  wire [64:0] _shiftReg_T_3 = enough ? _shiftReg_T_2 : hi; // @[src/main/scala/nutcore/backend/fu/MDU.scala 116:24]
  wire [128:0] _shiftReg_T_5 = {_shiftReg_T_3[63:0],lo,enough}; // @[src/main/scala/nutcore/backend/fu/MDU.scala 116:20]
  wire  wrap = cnt_value == 6'h3f; // @[src/main/scala/chisel3/util/Counter.scala 73:24]
  wire [5:0] _value_T_4 = cnt_value + 6'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire [2:0] _GEN_4 = wrap ? 3'h4 : state; // @[src/main/scala/nutcore/backend/fu/MDU.scala 118:{36,44} 77:22]
  wire [2:0] _GEN_5 = state == 3'h4 ? 3'h0 : state; // @[src/main/scala/nutcore/backend/fu/MDU.scala 119:36 120:11 77:22]
  wire [5:0] _GEN_7 = state == 3'h3 ? _value_T_4 : cnt_value; // @[src/main/scala/nutcore/backend/fu/MDU.scala 114:37 src/main/scala/chisel3/util/Counter.scala 77:15 61:40]
  wire [2:0] _GEN_8 = state == 3'h3 ? _GEN_4 : _GEN_5; // @[src/main/scala/nutcore/backend/fu/MDU.scala 114:37]
  wire [5:0] _GEN_11 = state == 3'h2 ? cnt_value : _GEN_7; // @[src/main/scala/nutcore/backend/fu/MDU.scala 111:35 src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [6:0] _GEN_12 = state == 3'h1 ? _value_T_2 : {{1'd0}, _GEN_11}; // @[src/main/scala/nutcore/backend/fu/MDU.scala 109:15 97:34]
  wire [6:0] _GEN_16 = newReq ? {{1'd0}, cnt_value} : _GEN_12; // @[src/main/scala/nutcore/backend/fu/MDU.scala 95:17 src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [63:0] r = hi[64:1]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 123:13]
  wire [63:0] _resQ_T_1 = 64'h0 - lo; // @[src/main/scala/nutcore/backend/fu/MDU.scala 124:28]
  wire [63:0] resQ = qSignReg ? _resQ_T_1 : lo; // @[src/main/scala/nutcore/backend/fu/MDU.scala 124:17]
  wire [63:0] _resR_T_1 = 64'h0 - r; // @[src/main/scala/nutcore/backend/fu/MDU.scala 125:28]
  wire [63:0] resR = aSignReg ? _resR_T_1 : r; // @[src/main/scala/nutcore/backend/fu/MDU.scala 125:17]
  wire [6:0] _GEN_21 = reset ? 7'h0 : _GEN_16; // @[src/main/scala/chisel3/util/Counter.scala 61:{40,40}]
  assign io_in_ready = state == 3'h0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 129:25]
  assign io_out_valid = state == 3'h4; // @[src/main/scala/nutcore/backend/fu/MDU.scala 128:39]
  assign io_out_bits = {resR,resQ}; // @[src/main/scala/nutcore/backend/fu/MDU.scala 126:21]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 77:22]
      state <= 3'h0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 77:22]
    end else if (newReq) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 95:17]
      state <= 3'h1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 96:11]
    end else if (state == 3'h1) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 97:34]
      state <= 3'h2; // @[src/main/scala/nutcore/backend/fu/MDU.scala 110:11]
    end else if (state == 3'h2) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 111:35]
      state <= 3'h3; // @[src/main/scala/nutcore/backend/fu/MDU.scala 113:11]
    end else begin
      state <= _GEN_8;
    end
    if (!(newReq)) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 95:17]
      if (!(state == 3'h1)) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 97:34]
        if (state == 3'h2) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 111:35]
          shiftReg <= {{1'd0}, _shiftReg_T}; // @[src/main/scala/nutcore/backend/fu/MDU.scala 112:14]
        end else if (state == 3'h3) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 114:37]
          shiftReg <= _shiftReg_T_5; // @[src/main/scala/nutcore/backend/fu/MDU.scala 116:14]
        end
      end
    end
    if (newReq) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 89:27]
      aSignReg <= aSign; // @[src/main/scala/nutcore/backend/fu/MDU.scala 89:27]
    end
    if (newReq) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 90:27]
      qSignReg <= (aSign ^ bSign) & ~divBy0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 90:27]
    end
    if (newReq) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
      if (bSign) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 73:12]
        bReg <= _T_3;
      end else begin
        bReg <= io_in_bits_1;
      end
    end
    if (newReq) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
      aValx2Reg <= _aValx2Reg_T; // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    cnt_value <= _GEN_21[5:0]; // @[src/main/scala/chisel3/util/Counter.scala 61:{40,40}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {5{`RANDOM}};
  shiftReg = _RAND_1[128:0];
  _RAND_2 = {1{`RANDOM}};
  aSignReg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  qSignReg = _RAND_3[0:0];
  _RAND_4 = {2{`RANDOM}};
  bReg = _RAND_4[63:0];
  _RAND_5 = {3{`RANDOM}};
  aValx2Reg = _RAND_5[64:0];
  _RAND_6 = {1{`RANDOM}};
  cnt_value = _RAND_6[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MDU(
  input         clock,
  input         reset,
  output        io_in_ready, // @[src/main/scala/nutcore/backend/fu/MDU.scala 136:14]
  input         io_in_valid, // @[src/main/scala/nutcore/backend/fu/MDU.scala 136:14]
  input  [63:0] io_in_bits_src1, // @[src/main/scala/nutcore/backend/fu/MDU.scala 136:14]
  input  [63:0] io_in_bits_src2, // @[src/main/scala/nutcore/backend/fu/MDU.scala 136:14]
  input  [6:0]  io_in_bits_func, // @[src/main/scala/nutcore/backend/fu/MDU.scala 136:14]
  input         io_out_ready, // @[src/main/scala/nutcore/backend/fu/MDU.scala 136:14]
  output        io_out_valid, // @[src/main/scala/nutcore/backend/fu/MDU.scala 136:14]
  output [63:0] io_out_bits // @[src/main/scala/nutcore/backend/fu/MDU.scala 136:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  mul_clock; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire  mul_reset; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire  mul_io_in_ready; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire  mul_io_in_valid; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire [64:0] mul_io_in_bits_0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire [64:0] mul_io_in_bits_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire  mul_io_out_ready; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire  mul_io_out_valid; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire [129:0] mul_io_out_bits; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire  div_clock; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire  div_reset; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire  div_io_in_ready; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire  div_io_in_valid; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire [63:0] div_io_in_bits_0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire [63:0] div_io_in_bits_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire  div_io_sign; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire  div_io_out_valid; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire [127:0] div_io_out_bits; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire  isDiv = io_in_bits_func[2]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 41:27]
  wire  isDivSign = isDiv & ~io_in_bits_func[0]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 42:39]
  wire  isW = io_in_bits_func[3]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 43:25]
  wire [64:0] _mul_io_in_bits_0_T_1 = {1'h0,io_in_bits_src1}; // @[src/main/scala/utils/BitUtils.scala 47:41]
  wire  mul_io_in_bits_0_signBit = io_in_bits_src1[63]; // @[src/main/scala/utils/BitUtils.scala 39:20]
  wire [64:0] _mul_io_in_bits_0_T_2 = {mul_io_in_bits_0_signBit,io_in_bits_src1}; // @[src/main/scala/utils/BitUtils.scala 40:41]
  wire  _mul_io_in_bits_0_T_5 = 2'h0 == io_in_bits_func[1:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _mul_io_in_bits_0_T_6 = 2'h1 == io_in_bits_func[1:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _mul_io_in_bits_0_T_7 = 2'h2 == io_in_bits_func[1:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _mul_io_in_bits_0_T_8 = 2'h3 == io_in_bits_func[1:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [64:0] _mul_io_in_bits_0_T_9 = _mul_io_in_bits_0_T_5 ? _mul_io_in_bits_0_T_1 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_0_T_10 = _mul_io_in_bits_0_T_6 ? _mul_io_in_bits_0_T_2 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_0_T_11 = _mul_io_in_bits_0_T_7 ? _mul_io_in_bits_0_T_2 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_0_T_12 = _mul_io_in_bits_0_T_8 ? _mul_io_in_bits_0_T_1 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_0_T_13 = _mul_io_in_bits_0_T_9 | _mul_io_in_bits_0_T_10; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_0_T_14 = _mul_io_in_bits_0_T_13 | _mul_io_in_bits_0_T_11; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_1_T_1 = {1'h0,io_in_bits_src2}; // @[src/main/scala/utils/BitUtils.scala 47:41]
  wire  mul_io_in_bits_1_signBit = io_in_bits_src2[63]; // @[src/main/scala/utils/BitUtils.scala 39:20]
  wire [64:0] _mul_io_in_bits_1_T_2 = {mul_io_in_bits_1_signBit,io_in_bits_src2}; // @[src/main/scala/utils/BitUtils.scala 40:41]
  wire [64:0] _mul_io_in_bits_1_T_9 = _mul_io_in_bits_0_T_5 ? _mul_io_in_bits_1_T_1 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_1_T_10 = _mul_io_in_bits_0_T_6 ? _mul_io_in_bits_1_T_2 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_1_T_11 = _mul_io_in_bits_0_T_7 ? _mul_io_in_bits_1_T_1 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_1_T_12 = _mul_io_in_bits_0_T_8 ? _mul_io_in_bits_1_T_1 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_1_T_13 = _mul_io_in_bits_1_T_9 | _mul_io_in_bits_1_T_10; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_1_T_14 = _mul_io_in_bits_1_T_13 | _mul_io_in_bits_1_T_11; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  div_io_in_bits_0_signBit = io_in_bits_src1[31]; // @[src/main/scala/utils/BitUtils.scala 39:20]
  wire [31:0] _div_io_in_bits_0_T_2 = div_io_in_bits_0_signBit ? 32'hffffffff : 32'h0; // @[src/main/scala/utils/BitUtils.scala 40:46]
  wire [63:0] _div_io_in_bits_0_T_3 = {_div_io_in_bits_0_T_2,io_in_bits_src1[31:0]}; // @[src/main/scala/utils/BitUtils.scala 40:41]
  wire [63:0] _div_io_in_bits_0_T_5 = {32'h0,io_in_bits_src1[31:0]}; // @[src/main/scala/utils/BitUtils.scala 47:41]
  wire [63:0] _div_io_in_bits_0_T_6 = isDivSign ? _div_io_in_bits_0_T_3 : _div_io_in_bits_0_T_5; // @[src/main/scala/nutcore/backend/fu/MDU.scala 169:47]
  wire  div_io_in_bits_1_signBit = io_in_bits_src2[31]; // @[src/main/scala/utils/BitUtils.scala 39:20]
  wire [31:0] _div_io_in_bits_1_T_2 = div_io_in_bits_1_signBit ? 32'hffffffff : 32'h0; // @[src/main/scala/utils/BitUtils.scala 40:46]
  wire [63:0] _div_io_in_bits_1_T_3 = {_div_io_in_bits_1_T_2,io_in_bits_src2[31:0]}; // @[src/main/scala/utils/BitUtils.scala 40:41]
  wire [63:0] _div_io_in_bits_1_T_5 = {32'h0,io_in_bits_src2[31:0]}; // @[src/main/scala/utils/BitUtils.scala 47:41]
  wire [63:0] _div_io_in_bits_1_T_6 = isDivSign ? _div_io_in_bits_1_T_3 : _div_io_in_bits_1_T_5; // @[src/main/scala/nutcore/backend/fu/MDU.scala 169:47]
  wire [63:0] mulRes = io_in_bits_func[1:0] == 2'h0 ? mul_io_out_bits[63:0] : mul_io_out_bits[127:64]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 176:19]
  wire [63:0] divRes = io_in_bits_func[1] ? div_io_out_bits[127:64] : div_io_out_bits[63:0]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 177:19]
  wire [63:0] res = isDiv ? divRes : mulRes; // @[src/main/scala/nutcore/backend/fu/MDU.scala 178:16]
  wire  io_out_bits_signBit = res[31]; // @[src/main/scala/utils/BitUtils.scala 39:20]
  wire [31:0] _io_out_bits_T_2 = io_out_bits_signBit ? 32'hffffffff : 32'h0; // @[src/main/scala/utils/BitUtils.scala 40:46]
  wire [63:0] _io_out_bits_T_3 = {_io_out_bits_T_2,res[31:0]}; // @[src/main/scala/utils/BitUtils.scala 40:41]
  wire  _isDivReg_T = io_in_ready & io_in_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  isDivReg_REG; // @[src/main/scala/nutcore/backend/fu/MDU.scala 181:48]
  wire  isDivReg = _isDivReg_T ? isDiv : isDivReg_REG; // @[src/main/scala/nutcore/backend/fu/MDU.scala 181:21]
  wire  _T_5 = mul_io_out_ready & mul_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  Multiplier mul ( // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
    .clock(mul_clock),
    .reset(mul_reset),
    .io_in_ready(mul_io_in_ready),
    .io_in_valid(mul_io_in_valid),
    .io_in_bits_0(mul_io_in_bits_0),
    .io_in_bits_1(mul_io_in_bits_1),
    .io_out_ready(mul_io_out_ready),
    .io_out_valid(mul_io_out_valid),
    .io_out_bits(mul_io_out_bits)
  );
  Divider div ( // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
    .clock(div_clock),
    .reset(div_reset),
    .io_in_ready(div_io_in_ready),
    .io_in_valid(div_io_in_valid),
    .io_in_bits_0(div_io_in_bits_0),
    .io_in_bits_1(div_io_in_bits_1),
    .io_sign(div_io_sign),
    .io_out_valid(div_io_out_valid),
    .io_out_bits(div_io_out_bits)
  );
  assign io_in_ready = isDiv ? div_io_in_ready : mul_io_in_ready; // @[src/main/scala/nutcore/backend/fu/MDU.scala 182:21]
  assign io_out_valid = isDivReg ? div_io_out_valid : mul_io_out_valid; // @[src/main/scala/nutcore/backend/fu/MDU.scala 183:22]
  assign io_out_bits = isW ? _io_out_bits_T_3 : res; // @[src/main/scala/nutcore/backend/fu/MDU.scala 179:21]
  assign mul_clock = clock;
  assign mul_reset = reset;
  assign mul_io_in_valid = io_in_valid & ~isDiv; // @[src/main/scala/nutcore/backend/fu/MDU.scala 173:34]
  assign mul_io_in_bits_0 = _mul_io_in_bits_0_T_14 | _mul_io_in_bits_0_T_12; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign mul_io_in_bits_1 = _mul_io_in_bits_1_T_14 | _mul_io_in_bits_1_T_12; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign mul_io_out_ready = 1'h1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 155:17]
  assign div_clock = clock;
  assign div_reset = reset;
  assign div_io_in_valid = io_in_valid & isDiv; // @[src/main/scala/nutcore/backend/fu/MDU.scala 174:34]
  assign div_io_in_bits_0 = isW ? _div_io_in_bits_0_T_6 : io_in_bits_src1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 169:38]
  assign div_io_in_bits_1 = isW ? _div_io_in_bits_1_T_6 : io_in_bits_src2; // @[src/main/scala/nutcore/backend/fu/MDU.scala 169:38]
  assign div_io_sign = isDiv & ~io_in_bits_func[0]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 42:39]
  always @(posedge clock) begin
    isDivReg_REG <= io_in_bits_func[2]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 41:27]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  isDivReg_REG = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CSR(
  input         clock,
  input         reset,
  input         io_in_valid, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input  [63:0] io_in_bits_src1, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input  [63:0] io_in_bits_src2, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input  [6:0]  io_in_bits_func, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input         io_out_ready, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  output        io_out_valid, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  output [63:0] io_out_bits, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input  [63:0] io_cfIn_instr, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input  [38:0] io_cfIn_pc, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input         io_cfIn_exceptionVec_1, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input         io_cfIn_exceptionVec_2, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input         io_cfIn_exceptionVec_4, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input         io_cfIn_exceptionVec_6, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input         io_cfIn_intrVec_0, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input         io_cfIn_intrVec_1, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input         io_cfIn_intrVec_2, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input         io_cfIn_intrVec_3, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input         io_cfIn_intrVec_4, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input         io_cfIn_intrVec_5, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input         io_cfIn_intrVec_6, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input         io_cfIn_intrVec_7, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input         io_cfIn_intrVec_8, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input         io_cfIn_intrVec_9, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input         io_cfIn_intrVec_10, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input         io_cfIn_intrVec_11, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  output [38:0] io_redirect_target, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  output        io_redirect_valid, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input         io_instrValid, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  output        io_wenFix, // @[src/main/scala/nutcore/backend/fu/CSR.scala 193:14]
  input         set_lr,
  input         perfCntCondMinstret,
  output        REG_1,
  input  [63:0] LSUADDR,
  output [11:0] intrVec_0,
  input  [63:0] set_lr_addr,
  input         perfCntCondMultiCommit,
  input         set_lr_val,
  output [63:0] lrAddr_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [31:0] _RAND_33;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] mtvec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 252:22]
  reg [63:0] mcounteren; // @[src/main/scala/nutcore/backend/fu/CSR.scala 253:27]
  reg [63:0] mcause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 254:23]
  reg [63:0] mtval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 255:22]
  reg [63:0] mepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 256:21]
  reg [63:0] mie; // @[src/main/scala/nutcore/backend/fu/CSR.scala 258:20]
  reg [63:0] mipReg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 260:24]
  wire  mip_s_u = mipReg[0]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 262:47]
  wire  mip_s_s = mipReg[1]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 262:47]
  wire  mip_s_h = mipReg[2]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 262:47]
  wire  mip_s_m = mipReg[3]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 262:47]
  wire  mip_t_u = mipReg[4]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 262:47]
  wire  mip_t_s = mipReg[5]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 262:47]
  wire  mip_t_h = mipReg[6]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 262:47]
  wire  mip_t_m = mipReg[7]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 262:47]
  wire  mip_e_u = mipReg[8]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 262:47]
  wire  mip_e_s = mipReg[9]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 262:47]
  wire  mip_e_h = mipReg[10]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 262:47]
  wire  mip_e_m = mipReg[11]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 262:47]
  reg [63:0] misa; // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:21]
  reg [63:0] mstatus; // @[src/main/scala/nutcore/backend/fu/CSR.scala 278:24]
  wire  mstatusStruct_ie_u = mstatus[0]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 300:39]
  wire  mstatusStruct_ie_s = mstatus[1]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 300:39]
  wire  mstatusStruct_ie_h = mstatus[2]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 300:39]
  wire  mstatusStruct_ie_m = mstatus[3]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 300:39]
  wire  mstatusStruct_pie_u = mstatus[4]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 300:39]
  wire  mstatusStruct_pie_s = mstatus[5]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 300:39]
  wire  mstatusStruct_pie_h = mstatus[6]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 300:39]
  wire  mstatusStruct_pie_m = mstatus[7]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 300:39]
  wire  mstatusStruct_spp = mstatus[8]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 300:39]
  wire [1:0] mstatusStruct_hpp = mstatus[10:9]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 300:39]
  wire [1:0] mstatusStruct_mpp = mstatus[12:11]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 300:39]
  wire [1:0] mstatusStruct_fs = mstatus[14:13]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 300:39]
  wire [1:0] mstatusStruct_xs = mstatus[16:15]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 300:39]
  wire  mstatusStruct_mprv = mstatus[17]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 300:39]
  wire  mstatusStruct_sum = mstatus[18]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 300:39]
  wire  mstatusStruct_mxr = mstatus[19]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 300:39]
  wire  mstatusStruct_tvm = mstatus[20]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 300:39]
  wire  mstatusStruct_tw = mstatus[21]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 300:39]
  wire  mstatusStruct_tsr = mstatus[22]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 300:39]
  wire [8:0] mstatusStruct_pad0 = mstatus[31:23]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 300:39]
  wire [1:0] mstatusStruct_uxl = mstatus[33:32]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 300:39]
  wire [1:0] mstatusStruct_sxl = mstatus[35:34]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 300:39]
  wire [26:0] mstatusStruct_pad1 = mstatus[62:36]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 300:39]
  wire  mstatusStruct_sd = mstatus[63]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 300:39]
  reg [63:0] medeleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 307:24]
  reg [63:0] mideleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 308:24]
  reg [63:0] mscratch; // @[src/main/scala/nutcore/backend/fu/CSR.scala 309:25]
  reg [63:0] pmpcfg0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 311:24]
  reg [63:0] pmpcfg1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 312:24]
  reg [63:0] pmpcfg2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 313:24]
  reg [63:0] pmpcfg3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 314:24]
  reg [63:0] pmpaddr0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 315:25]
  reg [63:0] pmpaddr1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 316:25]
  reg [63:0] pmpaddr2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 317:25]
  reg [63:0] pmpaddr3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:25]
  reg [63:0] stvec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 332:22]
  reg [63:0] satp; // @[src/main/scala/nutcore/backend/fu/CSR.scala 340:21]
  reg [63:0] sepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 341:21]
  reg [63:0] scause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 342:23]
  reg [63:0] stval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 343:22]
  reg [63:0] sscratch; // @[src/main/scala/nutcore/backend/fu/CSR.scala 344:25]
  reg [63:0] scounteren; // @[src/main/scala/nutcore/backend/fu/CSR.scala 345:27]
  reg  lr; // @[src/main/scala/nutcore/backend/fu/CSR.scala 358:19]
  reg [63:0] lrAddr; // @[src/main/scala/nutcore/backend/fu/CSR.scala 359:23]
  reg [1:0] priviledgeMode; // @[src/main/scala/nutcore/backend/fu/CSR.scala 372:31]
  reg [63:0] perfCnts_0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 377:47]
  reg [63:0] perfCnts_1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 377:47]
  reg [63:0] perfCnts_2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 377:47]
  wire [5:0] lo = {mip_t_s,mip_t_u,mip_s_m,mip_s_h,mip_s_s,mip_s_u}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 420:27]
  wire [11:0] _T_27 = {mip_e_m,mip_e_h,mip_e_s,mip_e_u,mip_t_m,mip_t_h,lo}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 420:27]
  wire [11:0] addr = io_in_bits_src2[11:0]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 460:18]
  wire [63:0] csri = {59'h0,io_cfIn_instr[19:15]}; // @[src/main/scala/utils/BitUtils.scala 47:41]
  wire  _rdata_T_37 = 12'hf12 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_38 = 12'h180 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_75 = _rdata_T_38 ? satp : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_39 = 12'h3b1 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_76 = _rdata_T_39 ? pmpaddr1 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_112 = _rdata_T_75 | _rdata_T_76; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_40 = 12'h3a2 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_77 = _rdata_T_40 ? pmpcfg2 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_113 = _rdata_T_112 | _rdata_T_77; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_41 = 12'h140 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_78 = _rdata_T_41 ? sscratch : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_114 = _rdata_T_113 | _rdata_T_78; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_42 = 12'h302 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_79 = _rdata_T_42 ? medeleg : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_115 = _rdata_T_114 | _rdata_T_79; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_43 = 12'h105 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_80 = _rdata_T_43 ? stvec : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_116 = _rdata_T_115 | _rdata_T_80; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_44 = 12'h141 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_81 = _rdata_T_44 ? sepc : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_117 = _rdata_T_116 | _rdata_T_81; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_45 = 12'h342 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_82 = _rdata_T_45 ? mcause : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_118 = _rdata_T_117 | _rdata_T_82; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_46 = 12'h306 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_83 = _rdata_T_46 ? mcounteren : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_119 = _rdata_T_118 | _rdata_T_83; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_47 = 12'hf11 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_48 = 12'h104 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_11 = mie & 64'h222; // @[src/main/scala/utils/RegMap.scala 48:84]
  wire [63:0] _rdata_T_85 = _rdata_T_48 ? _rdata_T_11 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_121 = _rdata_T_119 | _rdata_T_85; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_49 = 12'h144 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [11:0] _rdata_T_12 = _T_27 & 12'h222; // @[src/main/scala/utils/RegMap.scala 48:84]
  wire [11:0] _rdata_T_86 = _rdata_T_49 ? _rdata_T_12 : 12'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_78 = {{52'd0}, _rdata_T_86}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_122 = _rdata_T_121 | _GEN_78; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_50 = 12'h100 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_13 = mstatus & 64'h80000003000de122; // @[src/main/scala/utils/RegMap.scala 48:84]
  wire [63:0] _rdata_T_87 = _rdata_T_50 ? _rdata_T_13 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_123 = _rdata_T_122 | _rdata_T_87; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_51 = 12'h305 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_88 = _rdata_T_51 ? mtvec : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_124 = _rdata_T_123 | _rdata_T_88; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_52 = 12'h304 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_89 = _rdata_T_52 ? mie : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_125 = _rdata_T_124 | _rdata_T_89; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_53 = 12'hb01 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_90 = _rdata_T_53 ? perfCnts_1 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_126 = _rdata_T_125 | _rdata_T_90; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_54 = 12'h3b3 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_91 = _rdata_T_54 ? pmpaddr3 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_127 = _rdata_T_126 | _rdata_T_91; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_55 = 12'h143 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_92 = _rdata_T_55 ? stval : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_128 = _rdata_T_127 | _rdata_T_92; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_56 = 12'h301 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_93 = _rdata_T_56 ? misa : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_129 = _rdata_T_128 | _rdata_T_93; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_57 = 12'h300 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_94 = _rdata_T_57 ? mstatus : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_130 = _rdata_T_129 | _rdata_T_94; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_58 = 12'hb00 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_95 = _rdata_T_58 ? perfCnts_0 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_131 = _rdata_T_130 | _rdata_T_95; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_59 = 12'h3b0 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_96 = _rdata_T_59 ? pmpaddr0 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_132 = _rdata_T_131 | _rdata_T_96; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_60 = 12'h344 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_23 = {{52'd0}, _T_27}; // @[src/main/scala/utils/RegMap.scala 48:84]
  wire [63:0] _rdata_T_97 = _rdata_T_60 ? _rdata_T_23 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_133 = _rdata_T_132 | _rdata_T_97; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_61 = 12'hb02 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_98 = _rdata_T_61 ? perfCnts_2 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_134 = _rdata_T_133 | _rdata_T_98; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_62 = 12'h3a3 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_99 = _rdata_T_62 ? pmpcfg3 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_135 = _rdata_T_134 | _rdata_T_99; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_63 = 12'h303 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_100 = _rdata_T_63 ? mideleg : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_136 = _rdata_T_135 | _rdata_T_100; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_64 = 12'h3b2 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_101 = _rdata_T_64 ? pmpaddr2 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_137 = _rdata_T_136 | _rdata_T_101; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_65 = 12'hf13 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_66 = 12'h3a1 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_103 = _rdata_T_66 ? pmpcfg1 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_139 = _rdata_T_137 | _rdata_T_103; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_67 = 12'h340 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_104 = _rdata_T_67 ? mscratch : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_140 = _rdata_T_139 | _rdata_T_104; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_68 = 12'hf14 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_69 = 12'h341 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_106 = _rdata_T_69 ? mepc : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_142 = _rdata_T_140 | _rdata_T_106; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_70 = 12'h343 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_107 = _rdata_T_70 ? mtval : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_143 = _rdata_T_142 | _rdata_T_107; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_71 = 12'h106 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_108 = _rdata_T_71 ? scounteren : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_144 = _rdata_T_143 | _rdata_T_108; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_72 = 12'h3a0 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_109 = _rdata_T_72 ? pmpcfg0 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_145 = _rdata_T_144 | _rdata_T_109; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_73 = 12'h142 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_110 = _rdata_T_73 ? scause : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] rdata = _rdata_T_145 | _rdata_T_110; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T = rdata | io_in_bits_src1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 465:30]
  wire [63:0] _wdata_T_1 = ~io_in_bits_src1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 466:32]
  wire [63:0] _wdata_T_2 = rdata & _wdata_T_1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 466:30]
  wire [63:0] _wdata_T_3 = rdata | csri; // @[src/main/scala/nutcore/backend/fu/CSR.scala 468:30]
  wire [63:0] _wdata_T_4 = ~csri; // @[src/main/scala/nutcore/backend/fu/CSR.scala 469:32]
  wire [63:0] _wdata_T_5 = rdata & _wdata_T_4; // @[src/main/scala/nutcore/backend/fu/CSR.scala 469:30]
  wire  _wdata_T_6 = 7'h1 == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _wdata_T_7 = 7'h2 == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _wdata_T_8 = 7'h3 == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _wdata_T_9 = 7'h5 == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _wdata_T_10 = 7'h6 == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _wdata_T_11 = 7'h7 == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _wdata_T_12 = _wdata_T_6 ? io_in_bits_src1 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_13 = _wdata_T_7 ? _wdata_T : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_14 = _wdata_T_8 ? _wdata_T_2 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_15 = _wdata_T_9 ? csri : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_16 = _wdata_T_10 ? _wdata_T_3 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_17 = _wdata_T_11 ? _wdata_T_5 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_18 = _wdata_T_12 | _wdata_T_13; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_19 = _wdata_T_18 | _wdata_T_14; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_20 = _wdata_T_19 | _wdata_T_15; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_21 = _wdata_T_20 | _wdata_T_16; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] wdata = _wdata_T_21 | _wdata_T_17; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  satpLegalMode = wdata[63:60] == 4'h0 | wdata[63:60] == 4'h8; // @[src/main/scala/nutcore/backend/fu/CSR.scala 473:69]
  wire  wen = io_in_valid & io_in_bits_func != 7'h0 & (addr != 12'h180 | satpLegalMode); // @[src/main/scala/nutcore/backend/fu/CSR.scala 476:47]
  wire  isIllegalMode = priviledgeMode < addr[9:8]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 477:39]
  wire  justRead = (io_in_bits_func == 7'h2 | io_in_bits_func == 7'h6) & io_in_bits_src1 == 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 478:70]
  wire  isIllegalWrite = wen & addr[11:10] == 2'h3 & ~justRead; // @[src/main/scala/nutcore/backend/fu/CSR.scala 479:58]
  wire  isIllegalAccess = isIllegalMode | isIllegalWrite; // @[src/main/scala/nutcore/backend/fu/CSR.scala 480:39]
  wire  _T_72 = wen & ~isIllegalAccess; // @[src/main/scala/nutcore/backend/fu/CSR.scala 482:51]
  wire  _T_73 = addr == 12'h180; // @[src/main/scala/utils/RegMap.scala 50:65]
  wire  _T_81 = addr == 12'h302; // @[src/main/scala/utils/RegMap.scala 50:65]
  wire [63:0] _medeleg_T = wdata & 64'hbbff; // @[src/main/scala/utils/BitUtils.scala 32:13]
  wire [63:0] _medeleg_T_2 = medeleg & 64'h4400; // @[src/main/scala/utils/BitUtils.scala 32:36]
  wire [63:0] _medeleg_T_3 = _medeleg_T | _medeleg_T_2; // @[src/main/scala/utils/BitUtils.scala 32:25]
  wire [63:0] _GEN_8 = _T_72 & addr == 12'h141 ? wdata : sepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 341:21 src/main/scala/utils/RegMap.scala 50:{72,76}]
  wire [63:0] _GEN_9 = _T_72 & addr == 12'h342 ? wdata : mcause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 254:23 src/main/scala/utils/RegMap.scala 50:{72,76}]
  wire [63:0] _mie_T = wdata & 64'h222; // @[src/main/scala/utils/BitUtils.scala 32:13]
  wire [63:0] _mie_T_2 = mie & 64'h1dd; // @[src/main/scala/utils/BitUtils.scala 32:36]
  wire [63:0] _mie_T_3 = _mie_T | _mie_T_2; // @[src/main/scala/utils/BitUtils.scala 32:25]
  wire [63:0] _mstatus_T = wdata & 64'hc6122; // @[src/main/scala/utils/BitUtils.scala 32:13]
  wire [63:0] _mstatus_T_2 = mstatus & 64'h39edd; // @[src/main/scala/utils/BitUtils.scala 32:36]
  wire [63:0] _mstatus_T_3 = _mstatus_T | _mstatus_T_2; // @[src/main/scala/utils/BitUtils.scala 32:25]
  wire [1:0] mstatus_mstatusOld_fs = _mstatus_T_3[14:13]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 302:47]
  wire [63:0] mstatus_mstatusNew = {mstatus_mstatusOld_fs == 2'h3,_mstatus_T_3[62:0]}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 303:25]
  wire [63:0] _GEN_12 = _T_72 & addr == 12'h100 ? mstatus_mstatusNew : mstatus; // @[src/main/scala/nutcore/backend/fu/CSR.scala 278:24 src/main/scala/utils/RegMap.scala 50:{72,76}]
  wire [63:0] _GEN_17 = _T_72 & addr == 12'h143 ? wdata : stval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 343:22 src/main/scala/utils/RegMap.scala 50:{72,76}]
  wire [1:0] mstatus_mstatusOld_1_fs = wdata[14:13]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 302:47]
  wire [63:0] mstatus_mstatusNew_1 = {mstatus_mstatusOld_1_fs == 2'h3,wdata[62:0]}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 303:25]
  wire [63:0] _GEN_19 = _T_72 & addr == 12'h300 ? mstatus_mstatusNew_1 : _GEN_12; // @[src/main/scala/utils/RegMap.scala 50:{72,76}]
  wire [63:0] _mideleg_T_2 = mideleg & 64'h1dd; // @[src/main/scala/utils/BitUtils.scala 32:36]
  wire [63:0] _mideleg_T_3 = _mie_T | _mideleg_T_2; // @[src/main/scala/utils/BitUtils.scala 32:25]
  wire [63:0] _GEN_28 = _T_72 & addr == 12'h341 ? wdata : mepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 256:21 src/main/scala/utils/RegMap.scala 50:{72,76}]
  wire [63:0] _GEN_29 = _T_72 & addr == 12'h343 ? wdata : mtval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 255:22 src/main/scala/utils/RegMap.scala 50:{72,76}]
  wire [63:0] _GEN_32 = _T_72 & addr == 12'h142 ? wdata : scause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 342:23 src/main/scala/utils/RegMap.scala 50:{72,76}]
  wire  _isIllegalAddr_illegalAddr_T_1 = _rdata_T_37 ? 1'h0 : 1'h1; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_3 = _rdata_T_38 ? 1'h0 : _isIllegalAddr_illegalAddr_T_1; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_5 = _rdata_T_39 ? 1'h0 : _isIllegalAddr_illegalAddr_T_3; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_7 = _rdata_T_40 ? 1'h0 : _isIllegalAddr_illegalAddr_T_5; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_9 = _rdata_T_41 ? 1'h0 : _isIllegalAddr_illegalAddr_T_7; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_11 = _rdata_T_42 ? 1'h0 : _isIllegalAddr_illegalAddr_T_9; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_13 = _rdata_T_43 ? 1'h0 : _isIllegalAddr_illegalAddr_T_11; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_15 = _rdata_T_44 ? 1'h0 : _isIllegalAddr_illegalAddr_T_13; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_17 = _rdata_T_45 ? 1'h0 : _isIllegalAddr_illegalAddr_T_15; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_19 = _rdata_T_46 ? 1'h0 : _isIllegalAddr_illegalAddr_T_17; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_21 = _rdata_T_47 ? 1'h0 : _isIllegalAddr_illegalAddr_T_19; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_23 = _rdata_T_48 ? 1'h0 : _isIllegalAddr_illegalAddr_T_21; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_25 = _rdata_T_49 ? 1'h0 : _isIllegalAddr_illegalAddr_T_23; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_27 = _rdata_T_50 ? 1'h0 : _isIllegalAddr_illegalAddr_T_25; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_29 = _rdata_T_51 ? 1'h0 : _isIllegalAddr_illegalAddr_T_27; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_31 = _rdata_T_52 ? 1'h0 : _isIllegalAddr_illegalAddr_T_29; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_33 = _rdata_T_53 ? 1'h0 : _isIllegalAddr_illegalAddr_T_31; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_35 = _rdata_T_54 ? 1'h0 : _isIllegalAddr_illegalAddr_T_33; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_37 = _rdata_T_55 ? 1'h0 : _isIllegalAddr_illegalAddr_T_35; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_39 = _rdata_T_56 ? 1'h0 : _isIllegalAddr_illegalAddr_T_37; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_41 = _rdata_T_57 ? 1'h0 : _isIllegalAddr_illegalAddr_T_39; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_43 = _rdata_T_58 ? 1'h0 : _isIllegalAddr_illegalAddr_T_41; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_45 = _rdata_T_59 ? 1'h0 : _isIllegalAddr_illegalAddr_T_43; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_47 = _rdata_T_60 ? 1'h0 : _isIllegalAddr_illegalAddr_T_45; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_49 = _rdata_T_61 ? 1'h0 : _isIllegalAddr_illegalAddr_T_47; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_51 = _rdata_T_62 ? 1'h0 : _isIllegalAddr_illegalAddr_T_49; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_53 = _rdata_T_63 ? 1'h0 : _isIllegalAddr_illegalAddr_T_51; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_55 = _rdata_T_64 ? 1'h0 : _isIllegalAddr_illegalAddr_T_53; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_57 = _rdata_T_65 ? 1'h0 : _isIllegalAddr_illegalAddr_T_55; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_59 = _rdata_T_66 ? 1'h0 : _isIllegalAddr_illegalAddr_T_57; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_61 = _rdata_T_67 ? 1'h0 : _isIllegalAddr_illegalAddr_T_59; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_63 = _rdata_T_68 ? 1'h0 : _isIllegalAddr_illegalAddr_T_61; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_65 = _rdata_T_69 ? 1'h0 : _isIllegalAddr_illegalAddr_T_63; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_67 = _rdata_T_70 ? 1'h0 : _isIllegalAddr_illegalAddr_T_65; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_69 = _rdata_T_71 ? 1'h0 : _isIllegalAddr_illegalAddr_T_67; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_71 = _rdata_T_72 ? 1'h0 : _isIllegalAddr_illegalAddr_T_69; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  isIllegalAddr = _rdata_T_73 ? 1'h0 : _isIllegalAddr_illegalAddr_T_71; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  resetSatp = _T_73 & wen; // @[src/main/scala/nutcore/backend/fu/CSR.scala 484:35]
  wire [63:0] _mipReg_T_1 = wdata & 64'h77f; // @[src/main/scala/utils/BitUtils.scala 32:13]
  wire [63:0] _mipReg_T_3 = mipReg & 64'h80; // @[src/main/scala/utils/BitUtils.scala 32:36]
  wire [63:0] _mipReg_T_4 = _mipReg_T_1 | _mipReg_T_3; // @[src/main/scala/utils/BitUtils.scala 32:25]
  wire [63:0] _mipReg_T_7 = mipReg & 64'h1dd; // @[src/main/scala/utils/BitUtils.scala 32:36]
  wire [63:0] _mipReg_T_8 = _mie_T | _mipReg_T_7; // @[src/main/scala/utils/BitUtils.scala 32:25]
  wire  _isEbreak_T_1 = io_in_bits_func == 7'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 497:46]
  wire  isEbreak = addr == 12'h1 & io_in_bits_func == 7'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 497:38]
  wire  isEcall = addr == 12'h0 & _isEbreak_T_1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 498:36]
  wire  isMret = _T_81 & _isEbreak_T_1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 499:36]
  wire  isSret = addr == 12'h102 & _isEbreak_T_1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 500:36]
  wire  isUret = addr == 12'h2 & _isEbreak_T_1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 501:36]
  wire  tval_signBit_1 = io_cfIn_pc[38]; // @[src/main/scala/utils/BitUtils.scala 39:20]
  wire [24:0] _tval_T_8 = tval_signBit_1 ? 25'h1ffffff : 25'h0; // @[src/main/scala/utils/BitUtils.scala 40:46]
  wire [63:0] _tval_T_9 = {_tval_T_8,io_cfIn_pc}; // @[src/main/scala/utils/BitUtils.scala 40:41]
  wire  _T_154 = priviledgeMode == 2'h3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 569:25]
  wire  _T_163 = io_cfIn_exceptionVec_4 | io_cfIn_exceptionVec_6; // @[src/main/scala/nutcore/backend/fu/CSR.scala 577:30]
  wire [38:0] dmemAddrMisalignedAddr = LSUADDR[38:0]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 546:36 564:28]
  wire  mtval_signBit = dmemAddrMisalignedAddr[38]; // @[src/main/scala/utils/BitUtils.scala 39:20]
  wire [24:0] _mtval_T_5 = mtval_signBit ? 25'h1ffffff : 25'h0; // @[src/main/scala/utils/BitUtils.scala 40:46]
  wire [63:0] _mtval_T_6 = {_mtval_T_5,dmemAddrMisalignedAddr}; // @[src/main/scala/utils/BitUtils.scala 40:41]
  wire [63:0] _GEN_39 = _T_163 ? _mtval_T_6 : _GEN_29; // @[src/main/scala/nutcore/backend/fu/CSR.scala 578:3 579:11]
  wire [63:0] ideleg = mideleg & _rdata_T_23; // @[src/main/scala/nutcore/backend/fu/CSR.scala 603:26]
  wire  _intrVecEnable_0_T = priviledgeMode == 2'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 604:72]
  wire  _intrVecEnable_0_T_6 = priviledgeMode < 2'h3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 605:106]
  wire  _intrVecEnable_0_T_7 = _T_154 & mstatusStruct_ie_m | priviledgeMode < 2'h3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 605:87]
  wire  intrVecEnable_0 = ideleg[0] ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 :
    _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 604:51]
  wire  intrVecEnable_1 = ideleg[1] ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 :
    _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 604:51]
  wire  intrVecEnable_2 = ideleg[2] ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 :
    _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 604:51]
  wire  intrVecEnable_3 = ideleg[3] ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 :
    _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 604:51]
  wire  intrVecEnable_4 = ideleg[4] ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 :
    _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 604:51]
  wire  intrVecEnable_5 = ideleg[5] ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 :
    _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 604:51]
  wire  intrVecEnable_6 = ideleg[6] ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 :
    _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 604:51]
  wire  intrVecEnable_7 = ideleg[7] ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 :
    _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 604:51]
  wire  intrVecEnable_8 = ideleg[8] ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 :
    _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 604:51]
  wire  intrVecEnable_9 = ideleg[9] ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 :
    _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 604:51]
  wire  intrVecEnable_10 = ideleg[10] ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 :
    _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 604:51]
  wire  intrVecEnable_11 = ideleg[11] ? priviledgeMode == 2'h1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 :
    _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 604:51]
  wire [11:0] _intrVec_T_2 = mie[11:0] & _T_27; // @[src/main/scala/nutcore/backend/fu/CSR.scala 609:27]
  wire [5:0] intrVec_lo_1 = {intrVecEnable_5,intrVecEnable_4,intrVecEnable_3,intrVecEnable_2,intrVecEnable_1,
    intrVecEnable_0}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 609:65]
  wire [11:0] _intrVec_T_3 = {intrVecEnable_11,intrVecEnable_10,intrVecEnable_9,intrVecEnable_8,intrVecEnable_7,
    intrVecEnable_6,intrVec_lo_1}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 609:65]
  wire [11:0] intrVec = _intrVec_T_2 & _intrVec_T_3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 609:49]
  wire [2:0] _intrNO_T = io_cfIn_intrVec_4 ? 3'h4 : 3'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 613:69]
  wire [3:0] _intrNO_T_1 = io_cfIn_intrVec_8 ? 4'h8 : {{1'd0}, _intrNO_T}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 613:69]
  wire [3:0] _intrNO_T_2 = io_cfIn_intrVec_0 ? 4'h0 : _intrNO_T_1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 613:69]
  wire [3:0] _intrNO_T_3 = io_cfIn_intrVec_5 ? 4'h5 : _intrNO_T_2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 613:69]
  wire [3:0] _intrNO_T_4 = io_cfIn_intrVec_9 ? 4'h9 : _intrNO_T_3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 613:69]
  wire [3:0] _intrNO_T_5 = io_cfIn_intrVec_1 ? 4'h1 : _intrNO_T_4; // @[src/main/scala/nutcore/backend/fu/CSR.scala 613:69]
  wire [3:0] _intrNO_T_6 = io_cfIn_intrVec_7 ? 4'h7 : _intrNO_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 613:69]
  wire [3:0] _intrNO_T_7 = io_cfIn_intrVec_11 ? 4'hb : _intrNO_T_6; // @[src/main/scala/nutcore/backend/fu/CSR.scala 613:69]
  wire [3:0] intrNO = io_cfIn_intrVec_3 ? 4'h3 : _intrNO_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 613:69]
  wire [5:0] raiseIntr_lo = {io_cfIn_intrVec_5,io_cfIn_intrVec_4,io_cfIn_intrVec_3,io_cfIn_intrVec_2,io_cfIn_intrVec_1,
    io_cfIn_intrVec_0}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 615:35]
  wire [11:0] _raiseIntr_T = {io_cfIn_intrVec_11,io_cfIn_intrVec_10,io_cfIn_intrVec_9,io_cfIn_intrVec_8,
    io_cfIn_intrVec_7,io_cfIn_intrVec_6,raiseIntr_lo}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 615:35]
  wire  raiseIntr = |_raiseIntr_T; // @[src/main/scala/nutcore/backend/fu/CSR.scala 615:42]
  wire  csrExceptionVec_3 = io_in_valid & isEbreak; // @[src/main/scala/nutcore/backend/fu/CSR.scala 622:46]
  wire  csrExceptionVec_11 = _T_154 & io_in_valid & isEcall; // @[src/main/scala/nutcore/backend/fu/CSR.scala 623:70]
  wire  csrExceptionVec_9 = _intrVecEnable_0_T & io_in_valid & isEcall; // @[src/main/scala/nutcore/backend/fu/CSR.scala 624:70]
  wire  csrExceptionVec_8 = priviledgeMode == 2'h0 & io_in_valid & isEcall; // @[src/main/scala/nutcore/backend/fu/CSR.scala 625:70]
  wire  csrExceptionVec_2 = (isIllegalAddr | isIllegalAccess) & wen; // @[src/main/scala/nutcore/backend/fu/CSR.scala 626:71]
  wire [15:0] _raiseExceptionVec_T = {4'h0,csrExceptionVec_11,1'h0,csrExceptionVec_9,csrExceptionVec_8,4'h0,
    csrExceptionVec_3,csrExceptionVec_2,2'h0}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 630:43]
  wire [15:0] _raiseExceptionVec_T_1 = {8'h0,1'h0,io_cfIn_exceptionVec_6,1'h0,io_cfIn_exceptionVec_4,1'h0,
    io_cfIn_exceptionVec_2,io_cfIn_exceptionVec_1,1'h0}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 630:68]
  wire [15:0] raiseExceptionVec = _raiseExceptionVec_T | _raiseExceptionVec_T_1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 630:50]
  wire  raiseException = |raiseExceptionVec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 631:42]
  wire [2:0] _exceptionNO_T_1 = raiseExceptionVec[5] ? 3'h5 : 3'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 632:74]
  wire [2:0] _exceptionNO_T_3 = raiseExceptionVec[7] ? 3'h7 : _exceptionNO_T_1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 632:74]
  wire [3:0] _exceptionNO_T_5 = raiseExceptionVec[13] ? 4'hd : {{1'd0}, _exceptionNO_T_3}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 632:74]
  wire [3:0] _exceptionNO_T_7 = raiseExceptionVec[15] ? 4'hf : _exceptionNO_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 632:74]
  wire [3:0] _exceptionNO_T_9 = raiseExceptionVec[4] ? 4'h4 : _exceptionNO_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 632:74]
  wire [3:0] _exceptionNO_T_11 = raiseExceptionVec[6] ? 4'h6 : _exceptionNO_T_9; // @[src/main/scala/nutcore/backend/fu/CSR.scala 632:74]
  wire [3:0] _exceptionNO_T_13 = raiseExceptionVec[8] ? 4'h8 : _exceptionNO_T_11; // @[src/main/scala/nutcore/backend/fu/CSR.scala 632:74]
  wire [3:0] _exceptionNO_T_15 = raiseExceptionVec[9] ? 4'h9 : _exceptionNO_T_13; // @[src/main/scala/nutcore/backend/fu/CSR.scala 632:74]
  wire [3:0] _exceptionNO_T_17 = raiseExceptionVec[11] ? 4'hb : _exceptionNO_T_15; // @[src/main/scala/nutcore/backend/fu/CSR.scala 632:74]
  wire [3:0] _exceptionNO_T_19 = raiseExceptionVec[0] ? 4'h0 : _exceptionNO_T_17; // @[src/main/scala/nutcore/backend/fu/CSR.scala 632:74]
  wire [3:0] _exceptionNO_T_21 = raiseExceptionVec[2] ? 4'h2 : _exceptionNO_T_19; // @[src/main/scala/nutcore/backend/fu/CSR.scala 632:74]
  wire [3:0] _exceptionNO_T_23 = raiseExceptionVec[1] ? 4'h1 : _exceptionNO_T_21; // @[src/main/scala/nutcore/backend/fu/CSR.scala 632:74]
  wire [3:0] _exceptionNO_T_25 = raiseExceptionVec[12] ? 4'hc : _exceptionNO_T_23; // @[src/main/scala/nutcore/backend/fu/CSR.scala 632:74]
  wire [3:0] exceptionNO = raiseExceptionVec[3] ? 4'h3 : _exceptionNO_T_25; // @[src/main/scala/nutcore/backend/fu/CSR.scala 632:74]
  wire [63:0] _causeNO_T = {raiseIntr, 63'h0}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 635:28]
  wire [3:0] _causeNO_T_1 = raiseIntr ? intrNO : exceptionNO; // @[src/main/scala/nutcore/backend/fu/CSR.scala 635:46]
  wire [63:0] _GEN_80 = {{60'd0}, _causeNO_T_1}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 635:41]
  wire [63:0] causeNO = _causeNO_T | _GEN_80; // @[src/main/scala/nutcore/backend/fu/CSR.scala 635:41]
  wire  raiseExceptionIntr = (raiseException | raiseIntr) & io_instrValid; // @[src/main/scala/nutcore/backend/fu/CSR.scala 638:58]
  wire [38:0] _io_redirect_target_T_1 = io_cfIn_pc + 39'h4; // @[src/main/scala/nutcore/backend/fu/CSR.scala 643:51]
  wire [63:0] deleg = raiseIntr ? mideleg : medeleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 653:18]
  wire [63:0] _delegS_T_1 = deleg >> causeNO[3:0]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 655:22]
  wire  delegS = _delegS_T_1[0] & _intrVecEnable_0_T_6; // @[src/main/scala/nutcore/backend/fu/CSR.scala 655:38]
  wire [63:0] _trapTarget_T = delegS ? stvec : mtvec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 659:20]
  wire [38:0] trapTarget = _trapTarget_T[38:0]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 659:42]
  wire [38:0] _GEN_47 = io_in_valid & isSret ? sepc[38:0] : mepc[38:0]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 677:26 687:15]
  wire [38:0] retTarget = io_in_valid & isUret ? 39'h0 : _GEN_47; // @[src/main/scala/nutcore/backend/fu/CSR.scala 690:26 698:15]
  wire [38:0] _io_redirect_target_T_2 = raiseExceptionIntr ? trapTarget : retTarget; // @[src/main/scala/nutcore/backend/fu/CSR.scala 643:61]
  wire  tvalWen = ~_T_163 | raiseIntr; // @[src/main/scala/nutcore/backend/fu/CSR.scala 656:130]
  wire [5:0] mstatus_lo_lo = {mstatusStruct_pie_s,mstatusStruct_pie_u,mstatusStruct_pie_m,mstatusStruct_ie_h,
    mstatusStruct_ie_s,mstatusStruct_ie_u}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 672:27]
  wire [14:0] mstatus_lo = {mstatusStruct_fs,2'h0,mstatusStruct_hpp,mstatusStruct_spp,1'h1,mstatusStruct_pie_h,
    mstatus_lo_lo}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 672:27]
  wire [6:0] mstatus_hi_lo = {mstatusStruct_tw,mstatusStruct_tvm,mstatusStruct_mxr,mstatusStruct_sum,mstatusStruct_mprv,
    mstatusStruct_xs}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 672:27]
  wire [63:0] _mstatus_T_8 = {mstatusStruct_sd,mstatusStruct_pad1,mstatusStruct_sxl,mstatusStruct_uxl,mstatusStruct_pad0
    ,mstatusStruct_tsr,mstatus_hi_lo,mstatus_lo}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 672:27]
  wire [1:0] _GEN_40 = io_in_valid & isMret ? mstatusStruct_mpp : priviledgeMode; // @[src/main/scala/nutcore/backend/fu/CSR.scala 664:26 669:20 372:31]
  wire [63:0] _GEN_41 = io_in_valid & isMret ? _mstatus_T_8 : _GEN_19; // @[src/main/scala/nutcore/backend/fu/CSR.scala 664:26 672:13]
  wire [1:0] _priviledgeMode_T = {1'h0,mstatusStruct_spp}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 682:26]
  wire [5:0] mstatus_lo_lo_1 = {1'h1,mstatusStruct_pie_u,mstatusStruct_ie_m,mstatusStruct_ie_h,mstatusStruct_pie_s,
    mstatusStruct_ie_u}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 685:27]
  wire [14:0] mstatus_lo_1 = {mstatusStruct_fs,mstatusStruct_mpp,mstatusStruct_hpp,1'h0,mstatusStruct_pie_m,
    mstatusStruct_pie_h,mstatus_lo_lo_1}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 685:27]
  wire [63:0] _mstatus_T_9 = {mstatusStruct_sd,mstatusStruct_pad1,mstatusStruct_sxl,mstatusStruct_uxl,mstatusStruct_pad0
    ,mstatusStruct_tsr,mstatus_hi_lo,mstatus_lo_1}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 685:27]
  wire [5:0] mstatus_lo_lo_2 = {mstatusStruct_pie_s,1'h1,mstatusStruct_ie_m,mstatusStruct_ie_h,mstatusStruct_ie_s,
    mstatusStruct_pie_u}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 697:27]
  wire [14:0] mstatus_lo_2 = {mstatusStruct_fs,mstatusStruct_mpp,mstatusStruct_hpp,mstatusStruct_spp,mstatusStruct_pie_m
    ,mstatusStruct_pie_h,mstatus_lo_lo_2}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 697:27]
  wire [63:0] _mstatus_T_10 = {mstatusStruct_sd,mstatusStruct_pad1,mstatusStruct_sxl,mstatusStruct_uxl,
    mstatusStruct_pad0,mstatusStruct_tsr,mstatus_hi_lo,mstatus_lo_2}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 697:27]
  wire [1:0] _GEN_55 = delegS ? priviledgeMode : {{1'd0}, mstatusStruct_spp}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 705:19 708:22 703:30]
  wire  mstatusNew_3_pie_s = delegS ? mstatusStruct_ie_s : mstatusStruct_pie_s; // @[src/main/scala/nutcore/backend/fu/CSR.scala 705:19 709:24 703:30]
  wire  mstatusNew_3_ie_s = delegS ? 1'h0 : mstatusStruct_ie_s; // @[src/main/scala/nutcore/backend/fu/CSR.scala 705:19 710:23 703:30]
  wire [1:0] mstatusNew_3_mpp = delegS ? mstatusStruct_mpp : priviledgeMode; // @[src/main/scala/nutcore/backend/fu/CSR.scala 705:19 703:30 718:22]
  wire  mstatusNew_3_pie_m = delegS ? mstatusStruct_pie_m : mstatusStruct_ie_m; // @[src/main/scala/nutcore/backend/fu/CSR.scala 705:19 703:30 719:24]
  wire  mstatusNew_3_ie_m = delegS & mstatusStruct_ie_m; // @[src/main/scala/nutcore/backend/fu/CSR.scala 705:19 703:30 720:23]
  wire [5:0] mstatus_lo_lo_3 = {mstatusNew_3_pie_s,mstatusStruct_pie_u,mstatusNew_3_ie_m,mstatusStruct_ie_h,
    mstatusNew_3_ie_s,mstatusStruct_ie_u}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 732:27]
  wire  mstatusNew_3_spp = _GEN_55[0]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 703:30]
  wire [14:0] mstatus_lo_3 = {mstatusStruct_fs,mstatusNew_3_mpp,mstatusStruct_hpp,mstatusNew_3_spp,mstatusNew_3_pie_m,
    mstatusStruct_pie_h,mstatus_lo_lo_3}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 732:27]
  wire [63:0] _mstatus_T_11 = {mstatusStruct_sd,mstatusStruct_pad1,mstatusStruct_sxl,mstatusStruct_uxl,
    mstatusStruct_pad0,mstatusStruct_tsr,mstatus_hi_lo,mstatus_lo_3}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 732:27]
  wire [63:0] _perfCnts_0_T_5 = perfCnts_0 + 64'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 841:71]
  wire  _WIRE = 1'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 856:{33,33}]
  wire [63:0] _perfCnts_2_T_5 = perfCnts_2 + 64'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 841:71]
  wire [63:0] _perfCnts_2_T_7 = perfCnts_2 + 64'h2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 849:86]
  reg  REG; // @[src/main/scala/nutcore/backend/fu/CSR.scala 975:36]
  assign io_out_valid = io_in_valid; // @[src/main/scala/nutcore/backend/fu/CSR.scala 736:16]
  assign io_out_bits = _rdata_T_145 | _rdata_T_110; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_redirect_target = resetSatp ? _io_redirect_target_T_1 : _io_redirect_target_T_2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 643:28]
  assign io_redirect_valid = io_in_valid & _isEbreak_T_1 | raiseExceptionIntr | resetSatp; // @[src/main/scala/nutcore/backend/fu/CSR.scala 641:80]
  assign io_wenFix = |raiseExceptionVec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 631:42]
  assign REG_1 = REG;
  assign intrVec_0 = intrVec;
  assign lrAddr_0 = lrAddr;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 252:22]
      mtvec <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 252:22]
    end else if (_T_72 & addr == 12'h305) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      mtvec <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 253:27]
      mcounteren <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 253:27]
    end else if (_T_72 & addr == 12'h306) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      mcounteren <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 254:23]
      mcause <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 254:23]
    end else if (raiseExceptionIntr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 701:29]
      if (delegS) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 705:19]
        mcause <= _GEN_9;
      end else begin
        mcause <= causeNO; // @[src/main/scala/nutcore/backend/fu/CSR.scala 716:14]
      end
    end else begin
      mcause <= _GEN_9;
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 255:22]
      mtval <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 255:22]
    end else if (raiseExceptionIntr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 701:29]
      if (delegS) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 705:19]
        mtval <= _GEN_39;
      end else if (tvalWen) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 722:20]
        mtval <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 722:27]
      end else begin
        mtval <= _GEN_39;
      end
    end else begin
      mtval <= _GEN_39;
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 256:21]
      mepc <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 256:21]
    end else if (raiseExceptionIntr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 701:29]
      if (delegS) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 705:19]
        mepc <= _GEN_28;
      end else begin
        mepc <= _tval_T_9; // @[src/main/scala/nutcore/backend/fu/CSR.scala 717:12]
      end
    end else begin
      mepc <= _GEN_28;
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 258:20]
      mie <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 258:20]
    end else if (_T_72 & addr == 12'h304) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      mie <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end else if (_T_72 & addr == 12'h104) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      mie <= _mie_T_3; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 260:24]
      mipReg <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 260:24]
    end else if (_T_72 & addr == 12'h144) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      mipReg <= _mipReg_T_8; // @[src/main/scala/utils/RegMap.scala 50:76]
    end else if (_T_72 & addr == 12'h344) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      mipReg <= _mipReg_T_4; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:21]
      misa <= 64'h8000000000141101; // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:21]
    end else if (_T_72 & addr == 12'h301) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      misa <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 278:24]
      mstatus <= 64'h1800; // @[src/main/scala/nutcore/backend/fu/CSR.scala 278:24]
    end else if (raiseExceptionIntr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 701:29]
      mstatus <= _mstatus_T_11; // @[src/main/scala/nutcore/backend/fu/CSR.scala 732:13]
    end else if (io_in_valid & isUret) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 690:26]
      mstatus <= _mstatus_T_10; // @[src/main/scala/nutcore/backend/fu/CSR.scala 697:13]
    end else if (io_in_valid & isSret) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 677:26]
      mstatus <= _mstatus_T_9; // @[src/main/scala/nutcore/backend/fu/CSR.scala 685:13]
    end else begin
      mstatus <= _GEN_41;
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 307:24]
      medeleg <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 307:24]
    end else if (_T_72 & addr == 12'h302) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      medeleg <= _medeleg_T_3; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 308:24]
      mideleg <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 308:24]
    end else if (_T_72 & addr == 12'h303) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      mideleg <= _mideleg_T_3; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 309:25]
      mscratch <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 309:25]
    end else if (_T_72 & addr == 12'h340) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      mscratch <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 311:24]
      pmpcfg0 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 311:24]
    end else if (_T_72 & addr == 12'h3a0) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      pmpcfg0 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 312:24]
      pmpcfg1 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 312:24]
    end else if (_T_72 & addr == 12'h3a1) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      pmpcfg1 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 313:24]
      pmpcfg2 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 313:24]
    end else if (_T_72 & addr == 12'h3a2) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      pmpcfg2 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 314:24]
      pmpcfg3 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 314:24]
    end else if (_T_72 & addr == 12'h3a3) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      pmpcfg3 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 315:25]
      pmpaddr0 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 315:25]
    end else if (_T_72 & addr == 12'h3b0) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      pmpaddr0 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 316:25]
      pmpaddr1 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 316:25]
    end else if (_T_72 & addr == 12'h3b1) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      pmpaddr1 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 317:25]
      pmpaddr2 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 317:25]
    end else if (_T_72 & addr == 12'h3b2) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      pmpaddr2 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:25]
      pmpaddr3 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:25]
    end else if (_T_72 & addr == 12'h3b3) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      pmpaddr3 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 332:22]
      stvec <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 332:22]
    end else if (_T_72 & addr == 12'h105) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      stvec <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 340:21]
      satp <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 340:21]
    end else if (_T_72 & addr == 12'h180) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      satp <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 341:21]
      sepc <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 341:21]
    end else if (raiseExceptionIntr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 701:29]
      if (delegS) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 705:19]
        sepc <= _tval_T_9; // @[src/main/scala/nutcore/backend/fu/CSR.scala 707:12]
      end else begin
        sepc <= _GEN_8;
      end
    end else begin
      sepc <= _GEN_8;
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 342:23]
      scause <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 342:23]
    end else if (raiseExceptionIntr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 701:29]
      if (delegS) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 705:19]
        scause <= causeNO; // @[src/main/scala/nutcore/backend/fu/CSR.scala 706:14]
      end else begin
        scause <= _GEN_32;
      end
    end else begin
      scause <= _GEN_32;
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 343:22]
      stval <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 343:22]
    end else if (raiseExceptionIntr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 701:29]
      if (delegS) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 705:19]
        if (tvalWen) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 712:20]
          stval <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 712:27]
        end else begin
          stval <= _GEN_17;
        end
      end else begin
        stval <= _GEN_17;
      end
    end else begin
      stval <= _GEN_17;
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 344:25]
      sscratch <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 344:25]
    end else if (_T_72 & addr == 12'h140) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      sscratch <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 345:27]
      scounteren <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 345:27]
    end else if (_T_72 & addr == 12'h106) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      scounteren <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 358:19]
      lr <= 1'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 358:19]
    end else if (io_in_valid & isSret) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 677:26]
      lr <= 1'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 686:8]
    end else if (io_in_valid & isMret) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 664:26]
      lr <= 1'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 673:8]
    end else if (set_lr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 366:14]
      lr <= set_lr_val; // @[src/main/scala/nutcore/backend/fu/CSR.scala 367:8]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 359:23]
      lrAddr <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 359:23]
    end else if (set_lr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 366:14]
      lrAddr <= set_lr_addr; // @[src/main/scala/nutcore/backend/fu/CSR.scala 368:12]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 372:31]
      priviledgeMode <= 2'h3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 372:31]
    end else if (raiseExceptionIntr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 701:29]
      if (delegS) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 705:19]
        priviledgeMode <= 2'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 711:22]
      end else begin
        priviledgeMode <= 2'h3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 721:22]
      end
    end else if (io_in_valid & isUret) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 690:26]
      priviledgeMode <= 2'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 695:20]
    end else if (io_in_valid & isSret) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 677:26]
      priviledgeMode <= _priviledgeMode_T; // @[src/main/scala/nutcore/backend/fu/CSR.scala 682:20]
    end else begin
      priviledgeMode <= _GEN_40;
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 377:47]
      perfCnts_0 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 377:47]
    end else begin
      perfCnts_0 <= _perfCnts_0_T_5;
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 377:47]
      perfCnts_1 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 377:47]
    end else if (_T_72 & addr == 12'hb01) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_1 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 377:47]
      perfCnts_2 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 377:47]
    end else if (perfCntCondMultiCommit) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 849:35]
      perfCnts_2 <= _perfCnts_2_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 849:60]
    end else if (perfCntCondMinstret) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 841:62]
      perfCnts_2 <= _perfCnts_2_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 841:66]
    end else if (_T_72 & addr == 12'hb02) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_2 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 975:36]
      REG <= 1'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 975:36]
    end else begin
      REG <= raiseIntr & io_instrValid | raiseException & io_instrValid; // @[src/main/scala/nutcore/backend/fu/CSR.scala 975:36]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mtvec = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  mcounteren = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  mcause = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  mtval = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  mepc = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  mie = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  mipReg = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  misa = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  mstatus = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  medeleg = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  mideleg = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  mscratch = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  pmpcfg0 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  pmpcfg1 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  pmpcfg2 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  pmpcfg3 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  pmpaddr0 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  pmpaddr1 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  pmpaddr2 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  pmpaddr3 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  stvec = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  satp = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  sepc = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  scause = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  stval = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  sscratch = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  scounteren = _RAND_26[63:0];
  _RAND_27 = {1{`RANDOM}};
  lr = _RAND_27[0:0];
  _RAND_28 = {2{`RANDOM}};
  lrAddr = _RAND_28[63:0];
  _RAND_29 = {1{`RANDOM}};
  priviledgeMode = _RAND_29[1:0];
  _RAND_30 = {2{`RANDOM}};
  perfCnts_0 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  perfCnts_1 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  perfCnts_2 = _RAND_32[63:0];
  _RAND_33 = {1{`RANDOM}};
  REG = _RAND_33[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MOU(
  input         io_in_valid, // @[src/main/scala/nutcore/backend/fu/MOU.scala 38:14]
  input  [6:0]  io_in_bits_func, // @[src/main/scala/nutcore/backend/fu/MOU.scala 38:14]
  input  [38:0] io_cfIn_pc, // @[src/main/scala/nutcore/backend/fu/MOU.scala 38:14]
  output [38:0] io_redirect_target, // @[src/main/scala/nutcore/backend/fu/MOU.scala 38:14]
  output        io_redirect_valid, // @[src/main/scala/nutcore/backend/fu/MOU.scala 38:14]
  output        flushICache_0,
  output        flushTLB_0
);
  wire  flushICache = io_in_valid & io_in_bits_func == 7'h1; // @[src/main/scala/nutcore/backend/fu/MOU.scala 52:27]
  wire  flushTLB = io_in_valid & io_in_bits_func == 7'h2; // @[src/main/scala/nutcore/backend/fu/MOU.scala 56:24]
  assign io_redirect_target = io_cfIn_pc + 39'h4; // @[src/main/scala/nutcore/backend/fu/MOU.scala 49:36]
  assign io_redirect_valid = io_in_valid; // @[src/main/scala/nutcore/backend/fu/MOU.scala 50:21]
  assign flushICache_0 = flushICache;
  assign flushTLB_0 = flushTLB;
endmodule
module EXU(
  input         clock,
  input         reset,
  output        io_in_ready, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io_in_valid, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input  [63:0] io_in_bits_cf_instr, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input  [38:0] io_in_bits_cf_pc, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input  [38:0] io_in_bits_cf_pnpc, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io_in_bits_cf_exceptionVec_1, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io_in_bits_cf_exceptionVec_2, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io_in_bits_cf_intrVec_0, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io_in_bits_cf_intrVec_1, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io_in_bits_cf_intrVec_2, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io_in_bits_cf_intrVec_3, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io_in_bits_cf_intrVec_4, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io_in_bits_cf_intrVec_5, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io_in_bits_cf_intrVec_6, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io_in_bits_cf_intrVec_7, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io_in_bits_cf_intrVec_8, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io_in_bits_cf_intrVec_9, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io_in_bits_cf_intrVec_10, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io_in_bits_cf_intrVec_11, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input  [3:0]  io_in_bits_cf_brIdx, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input  [2:0]  io_in_bits_ctrl_fuType, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input  [6:0]  io_in_bits_ctrl_fuOpType, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input  [4:0]  io_in_bits_ctrl_rfSrc1, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input  [4:0]  io_in_bits_ctrl_rfSrc2, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io_in_bits_ctrl_rfWen, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input  [4:0]  io_in_bits_ctrl_rfDest, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input  [63:0] io_in_bits_data_src1, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input  [63:0] io_in_bits_data_src2, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input  [63:0] io_in_bits_data_imm, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io_out_ready, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output        io_out_valid, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [63:0] io_out_bits_decode_cf_instr, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [38:0] io_out_bits_decode_cf_pc, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [38:0] io_out_bits_decode_cf_redirect_target, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output        io_out_bits_decode_cf_redirect_valid, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [2:0]  io_out_bits_decode_ctrl_fuType, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [4:0]  io_out_bits_decode_ctrl_rfSrc1, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [4:0]  io_out_bits_decode_ctrl_rfSrc2, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output        io_out_bits_decode_ctrl_rfWen, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [4:0]  io_out_bits_decode_ctrl_rfDest, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [63:0] io_out_bits_decode_data_src1, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [63:0] io_out_bits_decode_data_src2, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [63:0] io_out_bits_commits_0, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [63:0] io_out_bits_commits_1, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [63:0] io_out_bits_commits_2, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [63:0] io_out_bits_commits_3, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [63:0] io_out_bits_mem_rvfi_addr_real, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [7:0]  io_out_bits_mem_rvfi_rmask, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [7:0]  io_out_bits_mem_rvfi_wmask, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [63:0] io_out_bits_mem_rvfi_rdata, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [63:0] io_out_bits_mem_rvfi_wdata, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io_flush, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io_dmem_req_ready, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output        io_dmem_req_valid, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [38:0] io_dmem_req_bits_addr, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [2:0]  io_dmem_req_bits_size, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [3:0]  io_dmem_req_bits_cmd, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [7:0]  io_dmem_req_bits_wmask, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [63:0] io_dmem_req_bits_wdata, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input         io_dmem_resp_valid, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  input  [63:0] io_dmem_resp_bits_rdata, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output        io_forward_valid, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output        io_forward_wb_rfWen, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [4:0]  io_forward_wb_rfDest, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [63:0] io_forward_wb_rfData, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output [2:0]  io_forward_fuType, // @[src/main/scala/nutcore/backend/seq/EXU.scala 29:14]
  output        _T_2_0,
  output        flushICache,
  output        REG_valid,
  output [38:0] REG_pc,
  output        REG_isMissPredict,
  output [38:0] REG_actualTarget,
  output        REG_actualTaken,
  output [6:0]  REG_fuOpType,
  output [1:0]  REG_btbType,
  output        REG_isRVC,
  input         io_in_valid_0,
  output        REG_0,
  output [11:0] intrVec,
  output        flushTLB,
  input         falseWire
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  alu_clock; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire  alu_reset; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire  alu_io_in_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire [63:0] alu_io_in_bits_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire [63:0] alu_io_in_bits_src2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire [6:0] alu_io_in_bits_func; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire  alu_io_out_ready; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire  alu_io_out_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire [63:0] alu_io_out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire [63:0] alu_io_cfIn_instr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire [38:0] alu_io_cfIn_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire [38:0] alu_io_cfIn_pnpc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire [3:0] alu_io_cfIn_brIdx; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire [38:0] alu_io_redirect_target; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire  alu_io_redirect_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire [63:0] alu_io_offset; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire  alu__T_2_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire  alu_REG_0_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire [38:0] alu_REG_0_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire  alu_REG_0_isMissPredict; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire [38:0] alu_REG_0_actualTarget; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire  alu_REG_0_actualTaken; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire [6:0] alu_REG_0_fuOpType; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire [1:0] alu_REG_0_btbType; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire  alu_REG_0_isRVC; // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
  wire  lsu_clock; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire  lsu_reset; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire  lsu_io__in_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire [63:0] lsu_io__in_bits_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire [63:0] lsu_io__in_bits_src2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire [6:0] lsu_io__in_bits_func; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire  lsu_io__out_ready; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire  lsu_io__out_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire [63:0] lsu_io__out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire [63:0] lsu_io__wdata; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire [31:0] lsu_io__instr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire  lsu_io__dmem_req_ready; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire  lsu_io__dmem_req_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire [38:0] lsu_io__dmem_req_bits_addr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire [2:0] lsu_io__dmem_req_bits_size; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire [3:0] lsu_io__dmem_req_bits_cmd; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire [7:0] lsu_io__dmem_req_bits_wmask; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire [63:0] lsu_io__dmem_req_bits_wdata; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire  lsu_io__dmem_resp_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire [63:0] lsu_io__dmem_resp_bits_rdata; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire  lsu_io__loadAddrMisaligned; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire  lsu_io__storeAddrMisaligned; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire  lsu_setLr_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire [63:0] lsu_io_in_bits_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire [63:0] lsu_setLrAddr_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire  lsu_setLrVal_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire [63:0] lsu_lr_addr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
  wire  mdu_clock; // @[src/main/scala/nutcore/backend/seq/EXU.scala 92:19]
  wire  mdu_reset; // @[src/main/scala/nutcore/backend/seq/EXU.scala 92:19]
  wire  mdu_io_in_ready; // @[src/main/scala/nutcore/backend/seq/EXU.scala 92:19]
  wire  mdu_io_in_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 92:19]
  wire [63:0] mdu_io_in_bits_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 92:19]
  wire [63:0] mdu_io_in_bits_src2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 92:19]
  wire [6:0] mdu_io_in_bits_func; // @[src/main/scala/nutcore/backend/seq/EXU.scala 92:19]
  wire  mdu_io_out_ready; // @[src/main/scala/nutcore/backend/seq/EXU.scala 92:19]
  wire  mdu_io_out_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 92:19]
  wire [63:0] mdu_io_out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 92:19]
  wire  csr_clock; // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:19]
  wire  csr_reset; // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:19]
  wire  csr_io_in_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:19]
  wire [63:0] csr_io_in_bits_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:19]
  wire [63:0] csr_io_in_bits_src2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:19]
  wire [6:0] csr_io_in_bits_func; // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:19]
  wire  csr_io_out_ready; // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:19]
  wire  csr_io_out_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:19]
  wire [63:0] csr_io_out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:19]
  wire [63:0] csr_io_cfIn_instr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:19]
  wire [38:0] csr_io_cfIn_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:19]
  wire  csr_io_cfIn_exceptionVec_1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:19]
  wire  csr_io_cfIn_exceptionVec_2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:19]
  wire  csr_io_cfIn_exceptionVec_4; // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:19]
  wire  csr_io_cfIn_exceptionVec_6; // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:19]
  wire  csr_io_cfIn_intrVec_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:19]
  wire  csr_io_cfIn_intrVec_1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:19]
  wire  csr_io_cfIn_intrVec_2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:19]
  wire  csr_io_cfIn_intrVec_3; // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:19]
  wire  csr_io_cfIn_intrVec_4; // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:19]
  wire  csr_io_cfIn_intrVec_5; // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:19]
  wire  csr_io_cfIn_intrVec_6; // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:19]
  wire  csr_io_cfIn_intrVec_7; // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:19]
  wire  csr_io_cfIn_intrVec_8; // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:19]
  wire  csr_io_cfIn_intrVec_9; // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:19]
  wire  csr_io_cfIn_intrVec_10; // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:19]
  wire  csr_io_cfIn_intrVec_11; // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:19]
  wire [38:0] csr_io_redirect_target; // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:19]
  wire  csr_io_redirect_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:19]
  wire  csr_io_instrValid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:19]
  wire  csr_io_wenFix; // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:19]
  wire  csr_set_lr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:19]
  wire  csr_perfCntCondMinstret; // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:19]
  wire  csr_REG_1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:19]
  wire [63:0] csr_LSUADDR; // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:19]
  wire [11:0] csr_intrVec_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:19]
  wire [63:0] csr_set_lr_addr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:19]
  wire  csr_perfCntCondMultiCommit; // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:19]
  wire  csr_set_lr_val; // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:19]
  wire [63:0] csr_lrAddr_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:19]
  wire  mou_io_in_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 111:19]
  wire [6:0] mou_io_in_bits_func; // @[src/main/scala/nutcore/backend/seq/EXU.scala 111:19]
  wire [38:0] mou_io_cfIn_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 111:19]
  wire [38:0] mou_io_redirect_target; // @[src/main/scala/nutcore/backend/seq/EXU.scala 111:19]
  wire  mou_io_redirect_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 111:19]
  wire  mou_flushICache_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 111:19]
  wire  mou_flushTLB_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 111:19]
  wire  _fuValids_0_T_2 = ~io_flush; // @[src/main/scala/nutcore/backend/seq/EXU.scala 44:84]
  wire  _fuValids_1_T = io_in_bits_ctrl_fuType == 3'h1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 44:57]
  wire  fuValids_1 = io_in_bits_ctrl_fuType == 3'h1 & io_in_valid & ~io_flush; // @[src/main/scala/nutcore/backend/seq/EXU.scala 44:81]
  wire  fuValids_3 = io_in_bits_ctrl_fuType == 3'h3 & io_in_valid & ~io_flush; // @[src/main/scala/nutcore/backend/seq/EXU.scala 44:81]
  reg [63:0] mem_rvfi_reg_addr_real; // @[src/main/scala/nutcore/backend/seq/EXU.scala 67:31]
  reg [7:0] mem_rvfi_reg_rmask; // @[src/main/scala/nutcore/backend/seq/EXU.scala 67:31]
  reg [7:0] mem_rvfi_reg_wmask; // @[src/main/scala/nutcore/backend/seq/EXU.scala 67:31]
  reg [63:0] mem_rvfi_reg_rdata; // @[src/main/scala/nutcore/backend/seq/EXU.scala 67:31]
  reg [63:0] mem_rvfi_reg_wdata; // @[src/main/scala/nutcore/backend/seq/EXU.scala 67:31]
  wire [7:0] _io_out_bits_mem_rvfi_rmask_T_1 = io_dmem_req_bits_cmd == 4'h0 ? io_dmem_req_bits_wmask : 8'h0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 73:42]
  wire [7:0] _io_out_bits_mem_rvfi_wmask_T_1 = io_dmem_req_bits_cmd == 4'h1 ? io_dmem_req_bits_wmask : 8'h0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 75:42]
  wire [63:0] _GEN_0 = io_dmem_req_valid ? {{25'd0}, io_dmem_req_bits_addr} : mem_rvfi_reg_addr_real; // @[src/main/scala/nutcore/backend/seq/EXU.scala 69:28 71:31 72:40]
  wire [7:0] _GEN_1 = io_dmem_req_valid ? _io_out_bits_mem_rvfi_rmask_T_1 : mem_rvfi_reg_rmask; // @[src/main/scala/nutcore/backend/seq/EXU.scala 69:28 71:31 73:36]
  wire [63:0] _GEN_2 = io_dmem_req_valid ? io_dmem_req_bits_wdata : mem_rvfi_reg_wdata; // @[src/main/scala/nutcore/backend/seq/EXU.scala 69:28 71:31 74:36]
  wire [7:0] _GEN_3 = io_dmem_req_valid ? _io_out_bits_mem_rvfi_wmask_T_1 : mem_rvfi_reg_wmask; // @[src/main/scala/nutcore/backend/seq/EXU.scala 69:28 71:31 75:36]
  wire [63:0] _GEN_6 = io_dmem_resp_valid ? io_dmem_resp_bits_rdata : mem_rvfi_reg_rdata; // @[src/main/scala/nutcore/backend/seq/EXU.scala 69:28 82:32 83:36]
  wire [38:0] _GEN_17 = csr_io_redirect_valid ? csr_io_redirect_target : alu_io_redirect_target; // @[src/main/scala/nutcore/backend/seq/EXU.scala 133:37 134:36 136:36]
  wire  _GEN_19 = csr_io_redirect_valid ? csr_io_redirect_valid : alu_io_redirect_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 133:37 134:36 136:36]
  wire  _io_out_valid_T_1 = 3'h1 == io_in_bits_ctrl_fuType ? lsu_io__out_valid : 1'h1; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _io_out_valid_T_3 = 3'h2 == io_in_bits_ctrl_fuType ? mdu_io_out_valid : _io_out_valid_T_1; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _io_forward_wb_rfData_T = alu_io_out_ready & alu_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  isBru = io_in_bits_ctrl_fuOpType[4]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 62:31]
  wire  _T_17 = _io_forward_wb_rfData_T & ~isBru; // @[src/main/scala/nutcore/backend/seq/EXU.scala 163:41]
  wire  _T_19 = _io_forward_wb_rfData_T & isBru; // @[src/main/scala/nutcore/backend/seq/EXU.scala 164:41]
  wire  _T_20 = lsu_io__out_ready & lsu_io__out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _T_21 = mdu_io_out_ready & mdu_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _T_22 = csr_io_out_ready & csr_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  ALU alu ( // @[src/main/scala/nutcore/backend/seq/EXU.scala 46:19]
    .clock(alu_clock),
    .reset(alu_reset),
    .io_in_valid(alu_io_in_valid),
    .io_in_bits_src1(alu_io_in_bits_src1),
    .io_in_bits_src2(alu_io_in_bits_src2),
    .io_in_bits_func(alu_io_in_bits_func),
    .io_out_ready(alu_io_out_ready),
    .io_out_valid(alu_io_out_valid),
    .io_out_bits(alu_io_out_bits),
    .io_cfIn_instr(alu_io_cfIn_instr),
    .io_cfIn_pc(alu_io_cfIn_pc),
    .io_cfIn_pnpc(alu_io_cfIn_pnpc),
    .io_cfIn_brIdx(alu_io_cfIn_brIdx),
    .io_redirect_target(alu_io_redirect_target),
    .io_redirect_valid(alu_io_redirect_valid),
    .io_offset(alu_io_offset),
    ._T_2_0(alu__T_2_0),
    .REG_0_valid(alu_REG_0_valid),
    .REG_0_pc(alu_REG_0_pc),
    .REG_0_isMissPredict(alu_REG_0_isMissPredict),
    .REG_0_actualTarget(alu_REG_0_actualTarget),
    .REG_0_actualTaken(alu_REG_0_actualTaken),
    .REG_0_fuOpType(alu_REG_0_fuOpType),
    .REG_0_btbType(alu_REG_0_btbType),
    .REG_0_isRVC(alu_REG_0_isRVC)
  );
  UnpipelinedLSU lsu ( // @[src/main/scala/nutcore/backend/seq/EXU.scala 54:19]
    .clock(lsu_clock),
    .reset(lsu_reset),
    .io__in_valid(lsu_io__in_valid),
    .io__in_bits_src1(lsu_io__in_bits_src1),
    .io__in_bits_src2(lsu_io__in_bits_src2),
    .io__in_bits_func(lsu_io__in_bits_func),
    .io__out_ready(lsu_io__out_ready),
    .io__out_valid(lsu_io__out_valid),
    .io__out_bits(lsu_io__out_bits),
    .io__wdata(lsu_io__wdata),
    .io__instr(lsu_io__instr),
    .io__dmem_req_ready(lsu_io__dmem_req_ready),
    .io__dmem_req_valid(lsu_io__dmem_req_valid),
    .io__dmem_req_bits_addr(lsu_io__dmem_req_bits_addr),
    .io__dmem_req_bits_size(lsu_io__dmem_req_bits_size),
    .io__dmem_req_bits_cmd(lsu_io__dmem_req_bits_cmd),
    .io__dmem_req_bits_wmask(lsu_io__dmem_req_bits_wmask),
    .io__dmem_req_bits_wdata(lsu_io__dmem_req_bits_wdata),
    .io__dmem_resp_valid(lsu_io__dmem_resp_valid),
    .io__dmem_resp_bits_rdata(lsu_io__dmem_resp_bits_rdata),
    .io__loadAddrMisaligned(lsu_io__loadAddrMisaligned),
    .io__storeAddrMisaligned(lsu_io__storeAddrMisaligned),
    .setLr_0(lsu_setLr_0),
    .io_in_bits_src1(lsu_io_in_bits_src1),
    .setLrAddr_0(lsu_setLrAddr_0),
    .setLrVal_0(lsu_setLrVal_0),
    .lr_addr(lsu_lr_addr)
  );
  MDU mdu ( // @[src/main/scala/nutcore/backend/seq/EXU.scala 92:19]
    .clock(mdu_clock),
    .reset(mdu_reset),
    .io_in_ready(mdu_io_in_ready),
    .io_in_valid(mdu_io_in_valid),
    .io_in_bits_src1(mdu_io_in_bits_src1),
    .io_in_bits_src2(mdu_io_in_bits_src2),
    .io_in_bits_func(mdu_io_in_bits_func),
    .io_out_ready(mdu_io_out_ready),
    .io_out_valid(mdu_io_out_valid),
    .io_out_bits(mdu_io_out_bits)
  );
  CSR csr ( // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:19]
    .clock(csr_clock),
    .reset(csr_reset),
    .io_in_valid(csr_io_in_valid),
    .io_in_bits_src1(csr_io_in_bits_src1),
    .io_in_bits_src2(csr_io_in_bits_src2),
    .io_in_bits_func(csr_io_in_bits_func),
    .io_out_ready(csr_io_out_ready),
    .io_out_valid(csr_io_out_valid),
    .io_out_bits(csr_io_out_bits),
    .io_cfIn_instr(csr_io_cfIn_instr),
    .io_cfIn_pc(csr_io_cfIn_pc),
    .io_cfIn_exceptionVec_1(csr_io_cfIn_exceptionVec_1),
    .io_cfIn_exceptionVec_2(csr_io_cfIn_exceptionVec_2),
    .io_cfIn_exceptionVec_4(csr_io_cfIn_exceptionVec_4),
    .io_cfIn_exceptionVec_6(csr_io_cfIn_exceptionVec_6),
    .io_cfIn_intrVec_0(csr_io_cfIn_intrVec_0),
    .io_cfIn_intrVec_1(csr_io_cfIn_intrVec_1),
    .io_cfIn_intrVec_2(csr_io_cfIn_intrVec_2),
    .io_cfIn_intrVec_3(csr_io_cfIn_intrVec_3),
    .io_cfIn_intrVec_4(csr_io_cfIn_intrVec_4),
    .io_cfIn_intrVec_5(csr_io_cfIn_intrVec_5),
    .io_cfIn_intrVec_6(csr_io_cfIn_intrVec_6),
    .io_cfIn_intrVec_7(csr_io_cfIn_intrVec_7),
    .io_cfIn_intrVec_8(csr_io_cfIn_intrVec_8),
    .io_cfIn_intrVec_9(csr_io_cfIn_intrVec_9),
    .io_cfIn_intrVec_10(csr_io_cfIn_intrVec_10),
    .io_cfIn_intrVec_11(csr_io_cfIn_intrVec_11),
    .io_redirect_target(csr_io_redirect_target),
    .io_redirect_valid(csr_io_redirect_valid),
    .io_instrValid(csr_io_instrValid),
    .io_wenFix(csr_io_wenFix),
    .set_lr(csr_set_lr),
    .perfCntCondMinstret(csr_perfCntCondMinstret),
    .REG_1(csr_REG_1),
    .LSUADDR(csr_LSUADDR),
    .intrVec_0(csr_intrVec_0),
    .set_lr_addr(csr_set_lr_addr),
    .perfCntCondMultiCommit(csr_perfCntCondMultiCommit),
    .set_lr_val(csr_set_lr_val),
    .lrAddr_0(csr_lrAddr_0)
  );
  MOU mou ( // @[src/main/scala/nutcore/backend/seq/EXU.scala 111:19]
    .io_in_valid(mou_io_in_valid),
    .io_in_bits_func(mou_io_in_bits_func),
    .io_cfIn_pc(mou_io_cfIn_pc),
    .io_redirect_target(mou_io_redirect_target),
    .io_redirect_valid(mou_io_redirect_valid),
    .flushICache_0(mou_flushICache_0),
    .flushTLB_0(mou_flushTLB_0)
  );
  assign io_in_ready = ~io_in_valid | io_out_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 154:31]
  assign io_out_valid = io_in_valid & _io_out_valid_T_3; // @[src/main/scala/nutcore/backend/seq/EXU.scala 143:31]
  assign io_out_bits_decode_cf_instr = io_in_bits_cf_instr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 128:31]
  assign io_out_bits_decode_cf_pc = io_in_bits_cf_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 127:28]
  assign io_out_bits_decode_cf_redirect_target = mou_io_redirect_valid ? mou_io_redirect_target : _GEN_17; // @[src/main/scala/nutcore/backend/seq/EXU.scala 131:32 132:36]
  assign io_out_bits_decode_cf_redirect_valid = mou_io_redirect_valid ? mou_io_redirect_valid : _GEN_19; // @[src/main/scala/nutcore/backend/seq/EXU.scala 131:32 132:36]
  assign io_out_bits_decode_ctrl_fuType = io_in_bits_ctrl_fuType; // @[src/main/scala/nutcore/backend/seq/EXU.scala 121:14]
  assign io_out_bits_decode_ctrl_rfSrc1 = io_in_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 122:14]
  assign io_out_bits_decode_ctrl_rfSrc2 = io_in_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 123:14]
  assign io_out_bits_decode_ctrl_rfWen = io_in_bits_ctrl_rfWen & (~lsu_io__loadAddrMisaligned & ~
    lsu_io__storeAddrMisaligned | ~fuValids_1) & ~(csr_io_wenFix & fuValids_3); // @[src/main/scala/nutcore/backend/seq/EXU.scala 119:125]
  assign io_out_bits_decode_ctrl_rfDest = io_in_bits_ctrl_rfDest; // @[src/main/scala/nutcore/backend/seq/EXU.scala 120:14]
  assign io_out_bits_decode_data_src1 = io_in_bits_ctrl_rfSrc1 == 5'h0 ? 64'h0 : io_in_bits_data_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 125:38]
  assign io_out_bits_decode_data_src2 = io_in_bits_ctrl_rfSrc2 == 5'h0 ? 64'h0 : io_in_bits_data_src2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 126:38]
  assign io_out_bits_commits_0 = alu_io_out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 148:35]
  assign io_out_bits_commits_1 = lsu_io__out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 149:35]
  assign io_out_bits_commits_2 = mdu_io_out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 151:35]
  assign io_out_bits_commits_3 = csr_io_out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 150:35]
  assign io_out_bits_mem_rvfi_addr_real = _fuValids_1_T ? _GEN_0 : 64'h0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:34 88:28]
  assign io_out_bits_mem_rvfi_rmask = _fuValids_1_T ? _GEN_1 : 8'h0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:34 88:28]
  assign io_out_bits_mem_rvfi_wmask = _fuValids_1_T ? _GEN_3 : 8'h0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:34 88:28]
  assign io_out_bits_mem_rvfi_rdata = _fuValids_1_T ? _GEN_6 : 64'h0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:34 88:28]
  assign io_out_bits_mem_rvfi_wdata = _fuValids_1_T ? _GEN_2 : 64'h0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:34 88:28]
  assign io_dmem_req_valid = lsu_io__dmem_req_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 60:11]
  assign io_dmem_req_bits_addr = lsu_io__dmem_req_bits_addr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 60:11]
  assign io_dmem_req_bits_size = lsu_io__dmem_req_bits_size; // @[src/main/scala/nutcore/backend/seq/EXU.scala 60:11]
  assign io_dmem_req_bits_cmd = lsu_io__dmem_req_bits_cmd; // @[src/main/scala/nutcore/backend/seq/EXU.scala 60:11]
  assign io_dmem_req_bits_wmask = lsu_io__dmem_req_bits_wmask; // @[src/main/scala/nutcore/backend/seq/EXU.scala 60:11]
  assign io_dmem_req_bits_wdata = lsu_io__dmem_req_bits_wdata; // @[src/main/scala/nutcore/backend/seq/EXU.scala 60:11]
  assign io_forward_valid = io_in_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 156:20]
  assign io_forward_wb_rfWen = io_in_bits_ctrl_rfWen; // @[src/main/scala/nutcore/backend/seq/EXU.scala 157:23]
  assign io_forward_wb_rfDest = io_in_bits_ctrl_rfDest; // @[src/main/scala/nutcore/backend/seq/EXU.scala 158:24]
  assign io_forward_wb_rfData = _io_forward_wb_rfData_T ? alu_io_out_bits : lsu_io__out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 159:30]
  assign io_forward_fuType = io_in_bits_ctrl_fuType; // @[src/main/scala/nutcore/backend/seq/EXU.scala 160:21]
  assign _T_2_0 = alu__T_2_0;
  assign flushICache = mou_flushICache_0;
  assign REG_valid = alu_REG_0_valid;
  assign REG_pc = alu_REG_0_pc;
  assign REG_isMissPredict = alu_REG_0_isMissPredict;
  assign REG_actualTarget = alu_REG_0_actualTarget;
  assign REG_actualTaken = alu_REG_0_actualTaken;
  assign REG_fuOpType = alu_REG_0_fuOpType;
  assign REG_btbType = alu_REG_0_btbType;
  assign REG_isRVC = alu_REG_0_isRVC;
  assign REG_0 = csr_REG_1;
  assign intrVec = csr_intrVec_0;
  assign flushTLB = mou_flushTLB_0;
  assign alu_clock = clock;
  assign alu_reset = reset;
  assign alu_io_in_valid = io_in_bits_ctrl_fuType == 3'h0 & io_in_valid & ~io_flush; // @[src/main/scala/nutcore/backend/seq/EXU.scala 44:81]
  assign alu_io_in_bits_src1 = io_in_bits_data_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 38:34]
  assign alu_io_in_bits_src2 = io_in_bits_data_src2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 39:34]
  assign alu_io_in_bits_func = io_in_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/fu/ALU.scala 83:15]
  assign alu_io_out_ready = 1'h1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 50:20]
  assign alu_io_cfIn_instr = io_in_bits_cf_instr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 48:15]
  assign alu_io_cfIn_pc = io_in_bits_cf_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 48:15]
  assign alu_io_cfIn_pnpc = io_in_bits_cf_pnpc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 48:15]
  assign alu_io_cfIn_brIdx = io_in_bits_cf_brIdx; // @[src/main/scala/nutcore/backend/seq/EXU.scala 48:15]
  assign alu_io_offset = io_in_bits_data_imm; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:17]
  assign lsu_clock = clock;
  assign lsu_reset = reset;
  assign lsu_io__in_valid = io_in_bits_ctrl_fuType == 3'h1 & io_in_valid & ~io_flush; // @[src/main/scala/nutcore/backend/seq/EXU.scala 44:81]
  assign lsu_io__in_bits_src1 = io_in_bits_data_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 38:34]
  assign lsu_io__in_bits_src2 = io_in_bits_data_imm; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 42:15]
  assign lsu_io__in_bits_func = io_in_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 43:15]
  assign lsu_io__out_ready = 1'h1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 61:20]
  assign lsu_io__wdata = io_in_bits_data_src2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 39:34]
  assign lsu_io__instr = io_in_bits_cf_instr[31:0]; // @[src/main/scala/nutcore/backend/seq/EXU.scala 58:16]
  assign lsu_io__dmem_req_ready = io_dmem_req_ready; // @[src/main/scala/nutcore/backend/seq/EXU.scala 60:11]
  assign lsu_io__dmem_resp_valid = io_dmem_resp_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 60:11]
  assign lsu_io__dmem_resp_bits_rdata = io_dmem_resp_bits_rdata; // @[src/main/scala/nutcore/backend/seq/EXU.scala 60:11]
  assign lsu_lr_addr = csr_lrAddr_0;
  assign mdu_clock = clock;
  assign mdu_reset = reset;
  assign mdu_io_in_valid = io_in_bits_ctrl_fuType == 3'h2 & io_in_valid & ~io_flush; // @[src/main/scala/nutcore/backend/seq/EXU.scala 44:81]
  assign mdu_io_in_bits_src1 = io_in_bits_data_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 38:34]
  assign mdu_io_in_bits_src2 = io_in_bits_data_src2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 39:34]
  assign mdu_io_in_bits_func = io_in_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/fu/MDU.scala 143:15]
  assign mdu_io_out_ready = 1'h1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 94:20]
  assign csr_clock = clock;
  assign csr_reset = reset;
  assign csr_io_in_valid = io_in_bits_ctrl_fuType == 3'h3 & io_in_valid & ~io_flush; // @[src/main/scala/nutcore/backend/seq/EXU.scala 44:81]
  assign csr_io_in_bits_src1 = io_in_bits_data_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 38:34]
  assign csr_io_in_bits_src2 = io_in_bits_data_src2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 39:34]
  assign csr_io_in_bits_func = io_in_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:15]
  assign csr_io_out_ready = 1'h1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 106:20]
  assign csr_io_cfIn_instr = io_in_bits_cf_instr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 99:15]
  assign csr_io_cfIn_pc = io_in_bits_cf_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 99:15]
  assign csr_io_cfIn_exceptionVec_1 = io_in_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 99:15]
  assign csr_io_cfIn_exceptionVec_2 = io_in_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 99:15]
  assign csr_io_cfIn_exceptionVec_4 = lsu_io__loadAddrMisaligned; // @[src/main/scala/nutcore/backend/seq/EXU.scala 100:48]
  assign csr_io_cfIn_exceptionVec_6 = lsu_io__storeAddrMisaligned; // @[src/main/scala/nutcore/backend/seq/EXU.scala 101:49]
  assign csr_io_cfIn_intrVec_0 = io_in_bits_cf_intrVec_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 99:15]
  assign csr_io_cfIn_intrVec_1 = io_in_bits_cf_intrVec_1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 99:15]
  assign csr_io_cfIn_intrVec_2 = io_in_bits_cf_intrVec_2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 99:15]
  assign csr_io_cfIn_intrVec_3 = io_in_bits_cf_intrVec_3; // @[src/main/scala/nutcore/backend/seq/EXU.scala 99:15]
  assign csr_io_cfIn_intrVec_4 = io_in_bits_cf_intrVec_4; // @[src/main/scala/nutcore/backend/seq/EXU.scala 99:15]
  assign csr_io_cfIn_intrVec_5 = io_in_bits_cf_intrVec_5; // @[src/main/scala/nutcore/backend/seq/EXU.scala 99:15]
  assign csr_io_cfIn_intrVec_6 = io_in_bits_cf_intrVec_6; // @[src/main/scala/nutcore/backend/seq/EXU.scala 99:15]
  assign csr_io_cfIn_intrVec_7 = io_in_bits_cf_intrVec_7; // @[src/main/scala/nutcore/backend/seq/EXU.scala 99:15]
  assign csr_io_cfIn_intrVec_8 = io_in_bits_cf_intrVec_8; // @[src/main/scala/nutcore/backend/seq/EXU.scala 99:15]
  assign csr_io_cfIn_intrVec_9 = io_in_bits_cf_intrVec_9; // @[src/main/scala/nutcore/backend/seq/EXU.scala 99:15]
  assign csr_io_cfIn_intrVec_10 = io_in_bits_cf_intrVec_10; // @[src/main/scala/nutcore/backend/seq/EXU.scala 99:15]
  assign csr_io_cfIn_intrVec_11 = io_in_bits_cf_intrVec_11; // @[src/main/scala/nutcore/backend/seq/EXU.scala 99:15]
  assign csr_io_instrValid = io_in_valid & _fuValids_0_T_2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 102:36]
  assign csr_set_lr = lsu_setLr_0;
  assign csr_perfCntCondMinstret = io_in_valid_0;
  assign csr_LSUADDR = lsu_io_in_bits_src1;
  assign csr_set_lr_addr = lsu_setLrAddr_0;
  assign csr_perfCntCondMultiCommit = falseWire;
  assign csr_set_lr_val = lsu_setLrVal_0;
  assign mou_io_in_valid = io_in_bits_ctrl_fuType == 3'h4 & io_in_valid & ~io_flush; // @[src/main/scala/nutcore/backend/seq/EXU.scala 44:81]
  assign mou_io_in_bits_func = io_in_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/fu/MOU.scala 45:15]
  assign mou_io_cfIn_pc = io_in_bits_cf_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 114:15]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/backend/seq/EXU.scala 67:31]
      mem_rvfi_reg_addr_real <= 64'h0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 67:31]
    end else if (_fuValids_1_T) begin // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:34]
      if (io_dmem_req_valid) begin // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:31]
        mem_rvfi_reg_addr_real <= {{25'd0}, io_dmem_req_bits_addr}; // @[src/main/scala/nutcore/backend/seq/EXU.scala 72:40]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/seq/EXU.scala 67:31]
      mem_rvfi_reg_rmask <= 8'h0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 67:31]
    end else if (_fuValids_1_T) begin // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:34]
      if (io_dmem_req_valid) begin // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:31]
        if (io_dmem_req_bits_cmd == 4'h0) begin // @[src/main/scala/nutcore/backend/seq/EXU.scala 73:42]
          mem_rvfi_reg_rmask <= io_dmem_req_bits_wmask;
        end else begin
          mem_rvfi_reg_rmask <= 8'h0;
        end
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/seq/EXU.scala 67:31]
      mem_rvfi_reg_wmask <= 8'h0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 67:31]
    end else if (_fuValids_1_T) begin // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:34]
      if (io_dmem_req_valid) begin // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:31]
        if (io_dmem_req_bits_cmd == 4'h1) begin // @[src/main/scala/nutcore/backend/seq/EXU.scala 75:42]
          mem_rvfi_reg_wmask <= io_dmem_req_bits_wmask;
        end else begin
          mem_rvfi_reg_wmask <= 8'h0;
        end
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/seq/EXU.scala 67:31]
      mem_rvfi_reg_rdata <= 64'h0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 67:31]
    end else if (_fuValids_1_T) begin // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:34]
      if (io_dmem_resp_valid) begin // @[src/main/scala/nutcore/backend/seq/EXU.scala 82:32]
        mem_rvfi_reg_rdata <= io_dmem_resp_bits_rdata; // @[src/main/scala/nutcore/backend/seq/EXU.scala 83:36]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/seq/EXU.scala 67:31]
      mem_rvfi_reg_wdata <= 64'h0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 67:31]
    end else if (_fuValids_1_T) begin // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:34]
      if (io_dmem_req_valid) begin // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:31]
        mem_rvfi_reg_wdata <= io_dmem_req_bits_wdata; // @[src/main/scala/nutcore/backend/seq/EXU.scala 74:36]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mem_rvfi_reg_addr_real = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  mem_rvfi_reg_rmask = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  mem_rvfi_reg_wmask = _RAND_2[7:0];
  _RAND_3 = {2{`RANDOM}};
  mem_rvfi_reg_rdata = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  mem_rvfi_reg_wdata = _RAND_4[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module WBU(
  input         clock,
  input         reset,
  input         io__in_valid, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [63:0] io__in_bits_decode_cf_instr, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [38:0] io__in_bits_decode_cf_pc, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [38:0] io__in_bits_decode_cf_redirect_target, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input         io__in_bits_decode_cf_redirect_valid, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [2:0]  io__in_bits_decode_ctrl_fuType, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [4:0]  io__in_bits_decode_ctrl_rfSrc1, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [4:0]  io__in_bits_decode_ctrl_rfSrc2, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input         io__in_bits_decode_ctrl_rfWen, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [4:0]  io__in_bits_decode_ctrl_rfDest, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [63:0] io__in_bits_decode_data_src1, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [63:0] io__in_bits_decode_data_src2, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [63:0] io__in_bits_commits_0, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [63:0] io__in_bits_commits_1, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [63:0] io__in_bits_commits_2, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [63:0] io__in_bits_commits_3, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [63:0] io__in_bits_mem_rvfi_addr_real, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [7:0]  io__in_bits_mem_rvfi_rmask, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [7:0]  io__in_bits_mem_rvfi_wmask, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [63:0] io__in_bits_mem_rvfi_rdata, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [63:0] io__in_bits_mem_rvfi_wdata, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  output        io__wb_rfWen, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  output [4:0]  io__wb_rfDest, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  output [63:0] io__wb_rfData, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  output [38:0] io__redirect_target, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  output        io__redirect_valid, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  output [63:0] io_in_bits_decode_data_src1,
  output        io_in_valid,
  output [4:0]  io_in_bits_decode_ctrl_rfSrc1,
  output [4:0]  io_wb_rfDest,
  output [63:0] rvfi_order_0,
  output [63:0] io_in_bits_mem_rvfi_addr_real,
  output [4:0]  io_in_bits_decode_ctrl_rfSrc2,
  output [63:0] _T_145_0,
  output        io_in_valid_0,
  output [63:0] io_in_bits_mem_rvfi_rdata,
  output [63:0] _T_151_0,
  output [63:0] io_in_bits_decode_cf_instr,
  output [63:0] io_in_bits_mem_rvfi_wdata,
  output [63:0] _T_142_0,
  output [63:0] io_in_bits_decode_data_src2,
  output [7:0]  io_in_bits_mem_rvfi_rmask,
  output        falseWire_0,
  output [7:0]  io_in_bits_mem_rvfi_wmask
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] _GEN_1 = 3'h1 == io__in_bits_decode_ctrl_fuType ? io__in_bits_commits_1 : io__in_bits_commits_0; // @[src/main/scala/nutcore/backend/seq/WBU.scala 37:{16,16}]
  wire [63:0] _GEN_2 = 3'h2 == io__in_bits_decode_ctrl_fuType ? io__in_bits_commits_2 : _GEN_1; // @[src/main/scala/nutcore/backend/seq/WBU.scala 37:{16,16}]
  wire [63:0] _GEN_3 = 3'h3 == io__in_bits_decode_ctrl_fuType ? io__in_bits_commits_3 : _GEN_2; // @[src/main/scala/nutcore/backend/seq/WBU.scala 37:{16,16}]
  wire  enableDisplay = 1'h0; // @[src/main/scala/utils/Debug.scala 40:{33,33}]
  wire [31:0] tmpInst = io__in_bits_decode_cf_instr[31:0]; // @[src/main/scala/nutcore/backend/seq/WBU.scala 104:47]
  wire [31:0] _T_6 = tmpInst & 32'h707f; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_7 = 32'h13 == _T_6; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_9 = 32'h2013 == _T_6; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_11 = 32'h3013 == _T_6; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_13 = 32'h7013 == _T_6; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_15 = 32'h6013 == _T_6; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_17 = 32'h4013 == _T_6; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [31:0] _T_18 = tmpInst & 32'hfc00707f; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 29:12]
  wire  _T_19 = 32'h1013 == _T_18; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 29:12]
  wire  _T_21 = 32'h5013 == _T_18; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 29:12]
  wire  _T_23 = 32'h40005013 == _T_18; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 29:12]
  wire [31:0] _T_24 = tmpInst & 32'h7f; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_25 = 32'h37 == _T_24; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_27 = 32'h17 == _T_24; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_29 = 32'h1b == _T_6; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire [31:0] _T_30 = tmpInst & 32'hfe00707f; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_31 = 32'h101b == _T_30; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_33 = 32'h501b == _T_30; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_37 = 32'h4000501b == _T_30; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_52 = _T_7 | _T_9 | _T_11 | _T_13 | _T_15 | _T_17 | _T_19 | _T_21 | _T_23 | _T_25 | _T_27 | _T_29 | _T_31 |
    _T_33 | _T_33 | _T_37; // @[riscv-spec-core/src/main/scala/rvspeccore/checker/AssumeHelper.scala 31:67]
  wire  _T_54 = 32'h33 == _T_30; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_56 = 32'h2033 == _T_30; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_58 = 32'h3033 == _T_30; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_60 = 32'h7033 == _T_30; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_62 = 32'h6033 == _T_30; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_64 = 32'h4033 == _T_30; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_66 = 32'h1033 == _T_30; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_68 = 32'h5033 == _T_30; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_70 = 32'h40000033 == _T_30; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_72 = 32'h40005033 == _T_30; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_81 = _T_54 | _T_56 | _T_58 | _T_60 | _T_62 | _T_64 | _T_66 | _T_68 | _T_70 | _T_72; // @[riscv-spec-core/src/main/scala/rvspeccore/checker/AssumeHelper.scala 31:67]
  wire  _T_84 = 32'h6f == _T_24; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_86 = 32'h67 == _T_6; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_88 = 32'h63 == _T_6; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_90 = 32'h1063 == _T_6; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_92 = 32'h4063 == _T_6; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_94 = 32'h6063 == _T_6; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_96 = 32'h5063 == _T_6; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_98 = 32'h7063 == _T_6; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_105 = _T_84 | _T_86 | _T_88 | _T_90 | _T_92 | _T_94 | _T_96 | _T_98; // @[riscv-spec-core/src/main/scala/rvspeccore/checker/AssumeHelper.scala 31:67]
  wire  _T_108 = 32'h3 == _T_6; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_110 = 32'h1003 == _T_6; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_112 = 32'h2003 == _T_6; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_114 = 32'h4003 == _T_6; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_116 = 32'h5003 == _T_6; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_118 = 32'h23 == _T_6; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_120 = 32'h1023 == _T_6; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_122 = 32'h2023 == _T_6; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_124 = 32'h6003 == _T_6; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_126 = 32'h3003 == _T_6; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_128 = 32'h3023 == _T_6; // @[riscv-spec-core/src/main/scala/rvspeccore/core/spec/RVInsts.scala 12:39]
  wire  _T_138 = _T_108 | _T_110 | _T_112 | _T_114 | _T_116 | _T_118 | _T_120 | _T_122 | _T_124 | _T_126 | _T_128; // @[riscv-spec-core/src/main/scala/rvspeccore/checker/AssumeHelper.scala 31:67]
  wire  _T_140 = ~io__in_valid | (_T_52 | _T_81 | _T_105 | _T_138); // @[src/main/scala/nutcore/backend/seq/WBU.scala 107:22]
  reg [63:0] rvfi_order; // @[src/main/scala/nutcore/backend/seq/WBU.scala 126:31]
  wire [63:0] _rvfi_order_T_1 = rvfi_order + 64'h1; // @[src/main/scala/nutcore/backend/seq/WBU.scala 128:34]
  wire [63:0] _T_142 = io__wb_rfDest == 5'h0 ? 64'h0 : io__wb_rfData; // @[src/main/scala/nutcore/backend/seq/WBU.scala 138:32]
  wire  signBit = io__in_bits_decode_cf_pc[38]; // @[src/main/scala/utils/BitUtils.scala 39:20]
  wire [24:0] _T_144 = signBit ? 25'h1ffffff : 25'h0; // @[src/main/scala/utils/BitUtils.scala 40:46]
  wire [63:0] _T_145 = {_T_144,io__in_bits_decode_cf_pc}; // @[src/main/scala/utils/BitUtils.scala 40:41]
  wire [63:0] _T_150 = _T_145 + 64'h4; // @[src/main/scala/nutcore/backend/seq/WBU.scala 141:95]
  wire [63:0] _T_151 = io__redirect_valid ? {{25'd0}, io__redirect_target} : _T_150; // @[src/main/scala/nutcore/backend/seq/WBU.scala 141:12]
  wire  falseWire = 1'h0; // @[src/main/scala/nutcore/backend/seq/WBU.scala 46:{27,27}]
  assign io__wb_rfWen = io__in_bits_decode_ctrl_rfWen & io__in_valid; // @[src/main/scala/nutcore/backend/seq/WBU.scala 35:47]
  assign io__wb_rfDest = io__in_bits_decode_ctrl_rfDest; // @[src/main/scala/nutcore/backend/seq/WBU.scala 36:16]
  assign io__wb_rfData = 3'h4 == io__in_bits_decode_ctrl_fuType ? 64'h0 : _GEN_3; // @[src/main/scala/nutcore/backend/seq/WBU.scala 37:{16,16}]
  assign io__redirect_target = io__in_bits_decode_cf_redirect_target; // @[src/main/scala/nutcore/backend/seq/WBU.scala 41:15]
  assign io__redirect_valid = io__in_bits_decode_cf_redirect_valid & io__in_valid; // @[src/main/scala/nutcore/backend/seq/WBU.scala 42:60]
  assign io_in_bits_decode_data_src1 = io__in_bits_decode_data_src1;
  assign io_in_valid = io__in_valid;
  assign io_in_bits_decode_ctrl_rfSrc1 = io__in_bits_decode_ctrl_rfSrc1;
  assign io_wb_rfDest = io__wb_rfDest;
  assign rvfi_order_0 = rvfi_order;
  assign io_in_bits_mem_rvfi_addr_real = io__in_bits_mem_rvfi_addr_real;
  assign io_in_bits_decode_ctrl_rfSrc2 = io__in_bits_decode_ctrl_rfSrc2;
  assign _T_145_0 = _T_145;
  assign io_in_valid_0 = io__in_valid;
  assign io_in_bits_mem_rvfi_rdata = io__in_bits_mem_rvfi_rdata;
  assign _T_151_0 = _T_151;
  assign io_in_bits_decode_cf_instr = io__in_bits_decode_cf_instr;
  assign io_in_bits_mem_rvfi_wdata = io__in_bits_mem_rvfi_wdata;
  assign _T_142_0 = _T_142;
  assign io_in_bits_decode_data_src2 = io__in_bits_decode_data_src2;
  assign io_in_bits_mem_rvfi_rmask = io__in_bits_mem_rvfi_rmask;
  assign falseWire_0 = enableDisplay;
  assign io_in_bits_mem_rvfi_wmask = io__in_bits_mem_rvfi_wmask;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/backend/seq/WBU.scala 126:31]
      rvfi_order <= 64'h0; // @[src/main/scala/nutcore/backend/seq/WBU.scala 126:31]
    end else if (io__in_valid) begin // @[src/main/scala/nutcore/backend/seq/WBU.scala 127:25]
      rvfi_order <= _rvfi_order_T_1; // @[src/main/scala/nutcore/backend/seq/WBU.scala 128:20]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  rvfi_order = _RAND_0[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Backend_inorder(
  input         clock,
  input         reset,
  output        io_in_0_ready, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 671:14]
  input         io_in_0_valid, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 671:14]
  input  [63:0] io_in_0_bits_cf_instr, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 671:14]
  input  [38:0] io_in_0_bits_cf_pc, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 671:14]
  input  [38:0] io_in_0_bits_cf_pnpc, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 671:14]
  input         io_in_0_bits_cf_exceptionVec_1, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 671:14]
  input         io_in_0_bits_cf_exceptionVec_2, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 671:14]
  input         io_in_0_bits_cf_intrVec_0, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 671:14]
  input         io_in_0_bits_cf_intrVec_1, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 671:14]
  input         io_in_0_bits_cf_intrVec_2, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 671:14]
  input         io_in_0_bits_cf_intrVec_3, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 671:14]
  input         io_in_0_bits_cf_intrVec_4, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 671:14]
  input         io_in_0_bits_cf_intrVec_5, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 671:14]
  input         io_in_0_bits_cf_intrVec_6, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 671:14]
  input         io_in_0_bits_cf_intrVec_7, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 671:14]
  input         io_in_0_bits_cf_intrVec_8, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 671:14]
  input         io_in_0_bits_cf_intrVec_9, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 671:14]
  input         io_in_0_bits_cf_intrVec_10, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 671:14]
  input         io_in_0_bits_cf_intrVec_11, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 671:14]
  input  [3:0]  io_in_0_bits_cf_brIdx, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 671:14]
  input         io_in_0_bits_ctrl_src1Type, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 671:14]
  input         io_in_0_bits_ctrl_src2Type, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 671:14]
  input  [2:0]  io_in_0_bits_ctrl_fuType, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 671:14]
  input  [6:0]  io_in_0_bits_ctrl_fuOpType, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 671:14]
  input  [4:0]  io_in_0_bits_ctrl_rfSrc1, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 671:14]
  input  [4:0]  io_in_0_bits_ctrl_rfSrc2, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 671:14]
  input         io_in_0_bits_ctrl_rfWen, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 671:14]
  input  [4:0]  io_in_0_bits_ctrl_rfDest, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 671:14]
  input  [63:0] io_in_0_bits_data_imm, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 671:14]
  input  [1:0]  io_flush, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 671:14]
  input         io_dmem_req_ready, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 671:14]
  output        io_dmem_req_valid, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 671:14]
  output [38:0] io_dmem_req_bits_addr, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 671:14]
  output [2:0]  io_dmem_req_bits_size, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 671:14]
  output [3:0]  io_dmem_req_bits_cmd, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 671:14]
  output [7:0]  io_dmem_req_bits_wmask, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 671:14]
  output [63:0] io_dmem_req_bits_wdata, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 671:14]
  input         io_dmem_resp_valid, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 671:14]
  input  [63:0] io_dmem_resp_bits_rdata, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 671:14]
  output [38:0] io_redirect_target, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 671:14]
  output        io_redirect_valid, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 671:14]
  output [63:0] io_in_bits_decode_data_src1,
  output        _T_2_0,
  output        io_in_valid,
  output [4:0]  io_in_bits_decode_ctrl_rfSrc1,
  output [4:0]  io_wb_rfDest,
  output        flushICache,
  output [63:0] rvfi_order,
  output [63:0] io_in_bits_mem_rvfi_addr_real,
  output [4:0]  io_in_bits_decode_ctrl_rfSrc2,
  output        REG_valid,
  output [38:0] REG_pc,
  output        REG_isMissPredict,
  output [38:0] REG_actualTarget,
  output        REG_actualTaken,
  output [6:0]  REG_fuOpType,
  output [1:0]  REG_btbType,
  output        REG_isRVC,
  output [63:0] _T_145,
  output [63:0] io_in_bits_mem_rvfi_rdata,
  output [63:0] _T_151,
  output [63:0] io_in_bits_decode_cf_instr,
  output        REG_0,
  output [63:0] io_in_bits_mem_rvfi_wdata,
  output [63:0] _T_142,
  output [63:0] io_in_bits_decode_data_src2,
  output [11:0] intrVec,
  output [7:0]  io_in_bits_mem_rvfi_rmask,
  output        flushTLB,
  output [7:0]  io_in_bits_mem_rvfi_wmask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
`endif // RANDOMIZE_REG_INIT
  wire  isu_clock; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  isu_reset; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  isu_io_in_0_ready; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  isu_io_in_0_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] isu_io_in_0_bits_cf_instr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [38:0] isu_io_in_0_bits_cf_pc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [38:0] isu_io_in_0_bits_cf_pnpc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  isu_io_in_0_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  isu_io_in_0_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  isu_io_in_0_bits_cf_intrVec_0; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  isu_io_in_0_bits_cf_intrVec_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  isu_io_in_0_bits_cf_intrVec_2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  isu_io_in_0_bits_cf_intrVec_3; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  isu_io_in_0_bits_cf_intrVec_4; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  isu_io_in_0_bits_cf_intrVec_5; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  isu_io_in_0_bits_cf_intrVec_6; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  isu_io_in_0_bits_cf_intrVec_7; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  isu_io_in_0_bits_cf_intrVec_8; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  isu_io_in_0_bits_cf_intrVec_9; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  isu_io_in_0_bits_cf_intrVec_10; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  isu_io_in_0_bits_cf_intrVec_11; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [3:0] isu_io_in_0_bits_cf_brIdx; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  isu_io_in_0_bits_ctrl_src1Type; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  isu_io_in_0_bits_ctrl_src2Type; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [2:0] isu_io_in_0_bits_ctrl_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [6:0] isu_io_in_0_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [4:0] isu_io_in_0_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [4:0] isu_io_in_0_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  isu_io_in_0_bits_ctrl_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [4:0] isu_io_in_0_bits_ctrl_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] isu_io_in_0_bits_data_imm; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  isu_io_out_ready; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  isu_io_out_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] isu_io_out_bits_cf_instr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [38:0] isu_io_out_bits_cf_pc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [38:0] isu_io_out_bits_cf_pnpc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  isu_io_out_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  isu_io_out_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  isu_io_out_bits_cf_intrVec_0; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  isu_io_out_bits_cf_intrVec_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  isu_io_out_bits_cf_intrVec_2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  isu_io_out_bits_cf_intrVec_3; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  isu_io_out_bits_cf_intrVec_4; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  isu_io_out_bits_cf_intrVec_5; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  isu_io_out_bits_cf_intrVec_6; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  isu_io_out_bits_cf_intrVec_7; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  isu_io_out_bits_cf_intrVec_8; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  isu_io_out_bits_cf_intrVec_9; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  isu_io_out_bits_cf_intrVec_10; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  isu_io_out_bits_cf_intrVec_11; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [3:0] isu_io_out_bits_cf_brIdx; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [2:0] isu_io_out_bits_ctrl_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [6:0] isu_io_out_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [4:0] isu_io_out_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [4:0] isu_io_out_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  isu_io_out_bits_ctrl_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [4:0] isu_io_out_bits_ctrl_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] isu_io_out_bits_data_src1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] isu_io_out_bits_data_src2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] isu_io_out_bits_data_imm; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  isu_io_wb_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [4:0] isu_io_wb_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] isu_io_wb_rfData; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  isu_io_forward_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  isu_io_forward_wb_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [4:0] isu_io_forward_wb_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] isu_io_forward_wb_rfData; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [2:0] isu_io_forward_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  isu_io_flush; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_clock; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  exu_reset; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  exu_io_in_ready; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  exu_io_in_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [63:0] exu_io_in_bits_cf_instr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [38:0] exu_io_in_bits_cf_pc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [38:0] exu_io_in_bits_cf_pnpc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  exu_io_in_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  exu_io_in_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  exu_io_in_bits_cf_intrVec_0; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  exu_io_in_bits_cf_intrVec_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  exu_io_in_bits_cf_intrVec_2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  exu_io_in_bits_cf_intrVec_3; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  exu_io_in_bits_cf_intrVec_4; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  exu_io_in_bits_cf_intrVec_5; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  exu_io_in_bits_cf_intrVec_6; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  exu_io_in_bits_cf_intrVec_7; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  exu_io_in_bits_cf_intrVec_8; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  exu_io_in_bits_cf_intrVec_9; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  exu_io_in_bits_cf_intrVec_10; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  exu_io_in_bits_cf_intrVec_11; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [3:0] exu_io_in_bits_cf_brIdx; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [2:0] exu_io_in_bits_ctrl_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [6:0] exu_io_in_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [4:0] exu_io_in_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [4:0] exu_io_in_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  exu_io_in_bits_ctrl_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [4:0] exu_io_in_bits_ctrl_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [63:0] exu_io_in_bits_data_src1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [63:0] exu_io_in_bits_data_src2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [63:0] exu_io_in_bits_data_imm; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  exu_io_out_ready; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  exu_io_out_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [63:0] exu_io_out_bits_decode_cf_instr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [38:0] exu_io_out_bits_decode_cf_pc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [38:0] exu_io_out_bits_decode_cf_redirect_target; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  exu_io_out_bits_decode_cf_redirect_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [2:0] exu_io_out_bits_decode_ctrl_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [4:0] exu_io_out_bits_decode_ctrl_rfSrc1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [4:0] exu_io_out_bits_decode_ctrl_rfSrc2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  exu_io_out_bits_decode_ctrl_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [4:0] exu_io_out_bits_decode_ctrl_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [63:0] exu_io_out_bits_decode_data_src1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [63:0] exu_io_out_bits_decode_data_src2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [63:0] exu_io_out_bits_commits_0; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [63:0] exu_io_out_bits_commits_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [63:0] exu_io_out_bits_commits_2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [63:0] exu_io_out_bits_commits_3; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [63:0] exu_io_out_bits_mem_rvfi_addr_real; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [7:0] exu_io_out_bits_mem_rvfi_rmask; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [7:0] exu_io_out_bits_mem_rvfi_wmask; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [63:0] exu_io_out_bits_mem_rvfi_rdata; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [63:0] exu_io_out_bits_mem_rvfi_wdata; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  exu_io_flush; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  exu_io_dmem_req_ready; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  exu_io_dmem_req_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [38:0] exu_io_dmem_req_bits_addr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [2:0] exu_io_dmem_req_bits_size; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [3:0] exu_io_dmem_req_bits_cmd; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [7:0] exu_io_dmem_req_bits_wmask; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [63:0] exu_io_dmem_req_bits_wdata; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  exu_io_dmem_resp_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [63:0] exu_io_dmem_resp_bits_rdata; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  exu_io_forward_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  exu_io_forward_wb_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [4:0] exu_io_forward_wb_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [63:0] exu_io_forward_wb_rfData; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [2:0] exu_io_forward_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  exu__T_2_0; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  exu_flushICache; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  exu_REG_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [38:0] exu_REG_pc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  exu_REG_isMissPredict; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [38:0] exu_REG_actualTarget; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  exu_REG_actualTaken; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [6:0] exu_REG_fuOpType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [1:0] exu_REG_btbType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  exu_REG_isRVC; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  exu_io_in_valid_0; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  exu_REG_0; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [11:0] exu_intrVec; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  exu_flushTLB; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  exu_falseWire; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  wbu_clock; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire  wbu_reset; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire  wbu_io__in_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire [63:0] wbu_io__in_bits_decode_cf_instr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire [38:0] wbu_io__in_bits_decode_cf_pc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire [38:0] wbu_io__in_bits_decode_cf_redirect_target; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire  wbu_io__in_bits_decode_cf_redirect_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire [2:0] wbu_io__in_bits_decode_ctrl_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire [4:0] wbu_io__in_bits_decode_ctrl_rfSrc1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire [4:0] wbu_io__in_bits_decode_ctrl_rfSrc2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire  wbu_io__in_bits_decode_ctrl_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire [4:0] wbu_io__in_bits_decode_ctrl_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire [63:0] wbu_io__in_bits_decode_data_src1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire [63:0] wbu_io__in_bits_decode_data_src2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire [63:0] wbu_io__in_bits_commits_0; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire [63:0] wbu_io__in_bits_commits_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire [63:0] wbu_io__in_bits_commits_2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire [63:0] wbu_io__in_bits_commits_3; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire [63:0] wbu_io__in_bits_mem_rvfi_addr_real; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire [7:0] wbu_io__in_bits_mem_rvfi_rmask; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire [7:0] wbu_io__in_bits_mem_rvfi_wmask; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire [63:0] wbu_io__in_bits_mem_rvfi_rdata; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire [63:0] wbu_io__in_bits_mem_rvfi_wdata; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire  wbu_io__wb_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire [4:0] wbu_io__wb_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire [63:0] wbu_io__wb_rfData; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire [38:0] wbu_io__redirect_target; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire  wbu_io__redirect_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire [63:0] wbu_io_in_bits_decode_data_src1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire  wbu_io_in_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire [4:0] wbu_io_in_bits_decode_ctrl_rfSrc1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire [4:0] wbu_io_wb_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire [63:0] wbu_rvfi_order_0; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire [63:0] wbu_io_in_bits_mem_rvfi_addr_real; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire [4:0] wbu_io_in_bits_decode_ctrl_rfSrc2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire [63:0] wbu__T_145_0; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire  wbu_io_in_valid_0; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire [63:0] wbu_io_in_bits_mem_rvfi_rdata; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire [63:0] wbu__T_151_0; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire [63:0] wbu_io_in_bits_decode_cf_instr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire [63:0] wbu_io_in_bits_mem_rvfi_wdata; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire [63:0] wbu__T_142_0; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire [63:0] wbu_io_in_bits_decode_data_src2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire [7:0] wbu_io_in_bits_mem_rvfi_rmask; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire  wbu_falseWire_0; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire [7:0] wbu_io_in_bits_mem_rvfi_wmask; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
  wire  _T = exu_io_out_ready & exu_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  valid; // @[src/main/scala/utils/Pipeline.scala 24:24]
  wire  _GEN_0 = _T ? 1'h0 : valid; // @[src/main/scala/utils/Pipeline.scala 24:24 25:{25,33}]
  wire  _T_2 = isu_io_out_valid & exu_io_in_ready; // @[src/main/scala/utils/Pipeline.scala 26:22]
  wire  _GEN_1 = isu_io_out_valid & exu_io_in_ready | _GEN_0; // @[src/main/scala/utils/Pipeline.scala 26:{38,46}]
  reg [63:0] exu_io_in_bits_r_cf_instr; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [38:0] exu_io_in_bits_r_cf_pc; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [38:0] exu_io_in_bits_r_cf_pnpc; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_exceptionVec_1; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_exceptionVec_2; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_intrVec_0; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_intrVec_1; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_intrVec_2; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_intrVec_3; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_intrVec_4; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_intrVec_5; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_intrVec_6; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_intrVec_7; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_intrVec_8; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_intrVec_9; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_intrVec_10; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_intrVec_11; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [3:0] exu_io_in_bits_r_cf_brIdx; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [2:0] exu_io_in_bits_r_ctrl_fuType; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [6:0] exu_io_in_bits_r_ctrl_fuOpType; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [4:0] exu_io_in_bits_r_ctrl_rfSrc1; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [4:0] exu_io_in_bits_r_ctrl_rfSrc2; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_ctrl_rfWen; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [4:0] exu_io_in_bits_r_ctrl_rfDest; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] exu_io_in_bits_r_data_src1; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] exu_io_in_bits_r_data_src2; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] exu_io_in_bits_r_data_imm; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  valid_1; // @[src/main/scala/utils/Pipeline.scala 24:24]
  wire  _T_4 = exu_io_out_valid; // @[src/main/scala/utils/Pipeline.scala 26:22]
  reg [63:0] wbu_io_in_bits_r_decode_cf_instr; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [38:0] wbu_io_in_bits_r_decode_cf_pc; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [38:0] wbu_io_in_bits_r_decode_cf_redirect_target; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  wbu_io_in_bits_r_decode_cf_redirect_valid; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [2:0] wbu_io_in_bits_r_decode_ctrl_fuType; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [4:0] wbu_io_in_bits_r_decode_ctrl_rfSrc1; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [4:0] wbu_io_in_bits_r_decode_ctrl_rfSrc2; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  wbu_io_in_bits_r_decode_ctrl_rfWen; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [4:0] wbu_io_in_bits_r_decode_ctrl_rfDest; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] wbu_io_in_bits_r_decode_data_src1; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] wbu_io_in_bits_r_decode_data_src2; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] wbu_io_in_bits_r_commits_0; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] wbu_io_in_bits_r_commits_1; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] wbu_io_in_bits_r_commits_2; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] wbu_io_in_bits_r_commits_3; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] wbu_io_in_bits_r_mem_rvfi_addr_real; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [7:0] wbu_io_in_bits_r_mem_rvfi_rmask; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [7:0] wbu_io_in_bits_r_mem_rvfi_wmask; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] wbu_io_in_bits_r_mem_rvfi_rdata; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] wbu_io_in_bits_r_mem_rvfi_wdata; // @[src/main/scala/utils/Pipeline.scala 30:28]
  ISU isu ( // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
    .clock(isu_clock),
    .reset(isu_reset),
    .io_in_0_ready(isu_io_in_0_ready),
    .io_in_0_valid(isu_io_in_0_valid),
    .io_in_0_bits_cf_instr(isu_io_in_0_bits_cf_instr),
    .io_in_0_bits_cf_pc(isu_io_in_0_bits_cf_pc),
    .io_in_0_bits_cf_pnpc(isu_io_in_0_bits_cf_pnpc),
    .io_in_0_bits_cf_exceptionVec_1(isu_io_in_0_bits_cf_exceptionVec_1),
    .io_in_0_bits_cf_exceptionVec_2(isu_io_in_0_bits_cf_exceptionVec_2),
    .io_in_0_bits_cf_intrVec_0(isu_io_in_0_bits_cf_intrVec_0),
    .io_in_0_bits_cf_intrVec_1(isu_io_in_0_bits_cf_intrVec_1),
    .io_in_0_bits_cf_intrVec_2(isu_io_in_0_bits_cf_intrVec_2),
    .io_in_0_bits_cf_intrVec_3(isu_io_in_0_bits_cf_intrVec_3),
    .io_in_0_bits_cf_intrVec_4(isu_io_in_0_bits_cf_intrVec_4),
    .io_in_0_bits_cf_intrVec_5(isu_io_in_0_bits_cf_intrVec_5),
    .io_in_0_bits_cf_intrVec_6(isu_io_in_0_bits_cf_intrVec_6),
    .io_in_0_bits_cf_intrVec_7(isu_io_in_0_bits_cf_intrVec_7),
    .io_in_0_bits_cf_intrVec_8(isu_io_in_0_bits_cf_intrVec_8),
    .io_in_0_bits_cf_intrVec_9(isu_io_in_0_bits_cf_intrVec_9),
    .io_in_0_bits_cf_intrVec_10(isu_io_in_0_bits_cf_intrVec_10),
    .io_in_0_bits_cf_intrVec_11(isu_io_in_0_bits_cf_intrVec_11),
    .io_in_0_bits_cf_brIdx(isu_io_in_0_bits_cf_brIdx),
    .io_in_0_bits_ctrl_src1Type(isu_io_in_0_bits_ctrl_src1Type),
    .io_in_0_bits_ctrl_src2Type(isu_io_in_0_bits_ctrl_src2Type),
    .io_in_0_bits_ctrl_fuType(isu_io_in_0_bits_ctrl_fuType),
    .io_in_0_bits_ctrl_fuOpType(isu_io_in_0_bits_ctrl_fuOpType),
    .io_in_0_bits_ctrl_rfSrc1(isu_io_in_0_bits_ctrl_rfSrc1),
    .io_in_0_bits_ctrl_rfSrc2(isu_io_in_0_bits_ctrl_rfSrc2),
    .io_in_0_bits_ctrl_rfWen(isu_io_in_0_bits_ctrl_rfWen),
    .io_in_0_bits_ctrl_rfDest(isu_io_in_0_bits_ctrl_rfDest),
    .io_in_0_bits_data_imm(isu_io_in_0_bits_data_imm),
    .io_out_ready(isu_io_out_ready),
    .io_out_valid(isu_io_out_valid),
    .io_out_bits_cf_instr(isu_io_out_bits_cf_instr),
    .io_out_bits_cf_pc(isu_io_out_bits_cf_pc),
    .io_out_bits_cf_pnpc(isu_io_out_bits_cf_pnpc),
    .io_out_bits_cf_exceptionVec_1(isu_io_out_bits_cf_exceptionVec_1),
    .io_out_bits_cf_exceptionVec_2(isu_io_out_bits_cf_exceptionVec_2),
    .io_out_bits_cf_intrVec_0(isu_io_out_bits_cf_intrVec_0),
    .io_out_bits_cf_intrVec_1(isu_io_out_bits_cf_intrVec_1),
    .io_out_bits_cf_intrVec_2(isu_io_out_bits_cf_intrVec_2),
    .io_out_bits_cf_intrVec_3(isu_io_out_bits_cf_intrVec_3),
    .io_out_bits_cf_intrVec_4(isu_io_out_bits_cf_intrVec_4),
    .io_out_bits_cf_intrVec_5(isu_io_out_bits_cf_intrVec_5),
    .io_out_bits_cf_intrVec_6(isu_io_out_bits_cf_intrVec_6),
    .io_out_bits_cf_intrVec_7(isu_io_out_bits_cf_intrVec_7),
    .io_out_bits_cf_intrVec_8(isu_io_out_bits_cf_intrVec_8),
    .io_out_bits_cf_intrVec_9(isu_io_out_bits_cf_intrVec_9),
    .io_out_bits_cf_intrVec_10(isu_io_out_bits_cf_intrVec_10),
    .io_out_bits_cf_intrVec_11(isu_io_out_bits_cf_intrVec_11),
    .io_out_bits_cf_brIdx(isu_io_out_bits_cf_brIdx),
    .io_out_bits_ctrl_fuType(isu_io_out_bits_ctrl_fuType),
    .io_out_bits_ctrl_fuOpType(isu_io_out_bits_ctrl_fuOpType),
    .io_out_bits_ctrl_rfSrc1(isu_io_out_bits_ctrl_rfSrc1),
    .io_out_bits_ctrl_rfSrc2(isu_io_out_bits_ctrl_rfSrc2),
    .io_out_bits_ctrl_rfWen(isu_io_out_bits_ctrl_rfWen),
    .io_out_bits_ctrl_rfDest(isu_io_out_bits_ctrl_rfDest),
    .io_out_bits_data_src1(isu_io_out_bits_data_src1),
    .io_out_bits_data_src2(isu_io_out_bits_data_src2),
    .io_out_bits_data_imm(isu_io_out_bits_data_imm),
    .io_wb_rfWen(isu_io_wb_rfWen),
    .io_wb_rfDest(isu_io_wb_rfDest),
    .io_wb_rfData(isu_io_wb_rfData),
    .io_forward_valid(isu_io_forward_valid),
    .io_forward_wb_rfWen(isu_io_forward_wb_rfWen),
    .io_forward_wb_rfDest(isu_io_forward_wb_rfDest),
    .io_forward_wb_rfData(isu_io_forward_wb_rfData),
    .io_forward_fuType(isu_io_forward_fuType),
    .io_flush(isu_io_flush)
  );
  EXU exu ( // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
    .clock(exu_clock),
    .reset(exu_reset),
    .io_in_ready(exu_io_in_ready),
    .io_in_valid(exu_io_in_valid),
    .io_in_bits_cf_instr(exu_io_in_bits_cf_instr),
    .io_in_bits_cf_pc(exu_io_in_bits_cf_pc),
    .io_in_bits_cf_pnpc(exu_io_in_bits_cf_pnpc),
    .io_in_bits_cf_exceptionVec_1(exu_io_in_bits_cf_exceptionVec_1),
    .io_in_bits_cf_exceptionVec_2(exu_io_in_bits_cf_exceptionVec_2),
    .io_in_bits_cf_intrVec_0(exu_io_in_bits_cf_intrVec_0),
    .io_in_bits_cf_intrVec_1(exu_io_in_bits_cf_intrVec_1),
    .io_in_bits_cf_intrVec_2(exu_io_in_bits_cf_intrVec_2),
    .io_in_bits_cf_intrVec_3(exu_io_in_bits_cf_intrVec_3),
    .io_in_bits_cf_intrVec_4(exu_io_in_bits_cf_intrVec_4),
    .io_in_bits_cf_intrVec_5(exu_io_in_bits_cf_intrVec_5),
    .io_in_bits_cf_intrVec_6(exu_io_in_bits_cf_intrVec_6),
    .io_in_bits_cf_intrVec_7(exu_io_in_bits_cf_intrVec_7),
    .io_in_bits_cf_intrVec_8(exu_io_in_bits_cf_intrVec_8),
    .io_in_bits_cf_intrVec_9(exu_io_in_bits_cf_intrVec_9),
    .io_in_bits_cf_intrVec_10(exu_io_in_bits_cf_intrVec_10),
    .io_in_bits_cf_intrVec_11(exu_io_in_bits_cf_intrVec_11),
    .io_in_bits_cf_brIdx(exu_io_in_bits_cf_brIdx),
    .io_in_bits_ctrl_fuType(exu_io_in_bits_ctrl_fuType),
    .io_in_bits_ctrl_fuOpType(exu_io_in_bits_ctrl_fuOpType),
    .io_in_bits_ctrl_rfSrc1(exu_io_in_bits_ctrl_rfSrc1),
    .io_in_bits_ctrl_rfSrc2(exu_io_in_bits_ctrl_rfSrc2),
    .io_in_bits_ctrl_rfWen(exu_io_in_bits_ctrl_rfWen),
    .io_in_bits_ctrl_rfDest(exu_io_in_bits_ctrl_rfDest),
    .io_in_bits_data_src1(exu_io_in_bits_data_src1),
    .io_in_bits_data_src2(exu_io_in_bits_data_src2),
    .io_in_bits_data_imm(exu_io_in_bits_data_imm),
    .io_out_ready(exu_io_out_ready),
    .io_out_valid(exu_io_out_valid),
    .io_out_bits_decode_cf_instr(exu_io_out_bits_decode_cf_instr),
    .io_out_bits_decode_cf_pc(exu_io_out_bits_decode_cf_pc),
    .io_out_bits_decode_cf_redirect_target(exu_io_out_bits_decode_cf_redirect_target),
    .io_out_bits_decode_cf_redirect_valid(exu_io_out_bits_decode_cf_redirect_valid),
    .io_out_bits_decode_ctrl_fuType(exu_io_out_bits_decode_ctrl_fuType),
    .io_out_bits_decode_ctrl_rfSrc1(exu_io_out_bits_decode_ctrl_rfSrc1),
    .io_out_bits_decode_ctrl_rfSrc2(exu_io_out_bits_decode_ctrl_rfSrc2),
    .io_out_bits_decode_ctrl_rfWen(exu_io_out_bits_decode_ctrl_rfWen),
    .io_out_bits_decode_ctrl_rfDest(exu_io_out_bits_decode_ctrl_rfDest),
    .io_out_bits_decode_data_src1(exu_io_out_bits_decode_data_src1),
    .io_out_bits_decode_data_src2(exu_io_out_bits_decode_data_src2),
    .io_out_bits_commits_0(exu_io_out_bits_commits_0),
    .io_out_bits_commits_1(exu_io_out_bits_commits_1),
    .io_out_bits_commits_2(exu_io_out_bits_commits_2),
    .io_out_bits_commits_3(exu_io_out_bits_commits_3),
    .io_out_bits_mem_rvfi_addr_real(exu_io_out_bits_mem_rvfi_addr_real),
    .io_out_bits_mem_rvfi_rmask(exu_io_out_bits_mem_rvfi_rmask),
    .io_out_bits_mem_rvfi_wmask(exu_io_out_bits_mem_rvfi_wmask),
    .io_out_bits_mem_rvfi_rdata(exu_io_out_bits_mem_rvfi_rdata),
    .io_out_bits_mem_rvfi_wdata(exu_io_out_bits_mem_rvfi_wdata),
    .io_flush(exu_io_flush),
    .io_dmem_req_ready(exu_io_dmem_req_ready),
    .io_dmem_req_valid(exu_io_dmem_req_valid),
    .io_dmem_req_bits_addr(exu_io_dmem_req_bits_addr),
    .io_dmem_req_bits_size(exu_io_dmem_req_bits_size),
    .io_dmem_req_bits_cmd(exu_io_dmem_req_bits_cmd),
    .io_dmem_req_bits_wmask(exu_io_dmem_req_bits_wmask),
    .io_dmem_req_bits_wdata(exu_io_dmem_req_bits_wdata),
    .io_dmem_resp_valid(exu_io_dmem_resp_valid),
    .io_dmem_resp_bits_rdata(exu_io_dmem_resp_bits_rdata),
    .io_forward_valid(exu_io_forward_valid),
    .io_forward_wb_rfWen(exu_io_forward_wb_rfWen),
    .io_forward_wb_rfDest(exu_io_forward_wb_rfDest),
    .io_forward_wb_rfData(exu_io_forward_wb_rfData),
    .io_forward_fuType(exu_io_forward_fuType),
    ._T_2_0(exu__T_2_0),
    .flushICache(exu_flushICache),
    .REG_valid(exu_REG_valid),
    .REG_pc(exu_REG_pc),
    .REG_isMissPredict(exu_REG_isMissPredict),
    .REG_actualTarget(exu_REG_actualTarget),
    .REG_actualTaken(exu_REG_actualTaken),
    .REG_fuOpType(exu_REG_fuOpType),
    .REG_btbType(exu_REG_btbType),
    .REG_isRVC(exu_REG_isRVC),
    .io_in_valid_0(exu_io_in_valid_0),
    .REG_0(exu_REG_0),
    .intrVec(exu_intrVec),
    .flushTLB(exu_flushTLB),
    .falseWire(exu_falseWire)
  );
  WBU wbu ( // @[src/main/scala/nutcore/backend/ooo/Backend.scala 682:20]
    .clock(wbu_clock),
    .reset(wbu_reset),
    .io__in_valid(wbu_io__in_valid),
    .io__in_bits_decode_cf_instr(wbu_io__in_bits_decode_cf_instr),
    .io__in_bits_decode_cf_pc(wbu_io__in_bits_decode_cf_pc),
    .io__in_bits_decode_cf_redirect_target(wbu_io__in_bits_decode_cf_redirect_target),
    .io__in_bits_decode_cf_redirect_valid(wbu_io__in_bits_decode_cf_redirect_valid),
    .io__in_bits_decode_ctrl_fuType(wbu_io__in_bits_decode_ctrl_fuType),
    .io__in_bits_decode_ctrl_rfSrc1(wbu_io__in_bits_decode_ctrl_rfSrc1),
    .io__in_bits_decode_ctrl_rfSrc2(wbu_io__in_bits_decode_ctrl_rfSrc2),
    .io__in_bits_decode_ctrl_rfWen(wbu_io__in_bits_decode_ctrl_rfWen),
    .io__in_bits_decode_ctrl_rfDest(wbu_io__in_bits_decode_ctrl_rfDest),
    .io__in_bits_decode_data_src1(wbu_io__in_bits_decode_data_src1),
    .io__in_bits_decode_data_src2(wbu_io__in_bits_decode_data_src2),
    .io__in_bits_commits_0(wbu_io__in_bits_commits_0),
    .io__in_bits_commits_1(wbu_io__in_bits_commits_1),
    .io__in_bits_commits_2(wbu_io__in_bits_commits_2),
    .io__in_bits_commits_3(wbu_io__in_bits_commits_3),
    .io__in_bits_mem_rvfi_addr_real(wbu_io__in_bits_mem_rvfi_addr_real),
    .io__in_bits_mem_rvfi_rmask(wbu_io__in_bits_mem_rvfi_rmask),
    .io__in_bits_mem_rvfi_wmask(wbu_io__in_bits_mem_rvfi_wmask),
    .io__in_bits_mem_rvfi_rdata(wbu_io__in_bits_mem_rvfi_rdata),
    .io__in_bits_mem_rvfi_wdata(wbu_io__in_bits_mem_rvfi_wdata),
    .io__wb_rfWen(wbu_io__wb_rfWen),
    .io__wb_rfDest(wbu_io__wb_rfDest),
    .io__wb_rfData(wbu_io__wb_rfData),
    .io__redirect_target(wbu_io__redirect_target),
    .io__redirect_valid(wbu_io__redirect_valid),
    .io_in_bits_decode_data_src1(wbu_io_in_bits_decode_data_src1),
    .io_in_valid(wbu_io_in_valid),
    .io_in_bits_decode_ctrl_rfSrc1(wbu_io_in_bits_decode_ctrl_rfSrc1),
    .io_wb_rfDest(wbu_io_wb_rfDest),
    .rvfi_order_0(wbu_rvfi_order_0),
    .io_in_bits_mem_rvfi_addr_real(wbu_io_in_bits_mem_rvfi_addr_real),
    .io_in_bits_decode_ctrl_rfSrc2(wbu_io_in_bits_decode_ctrl_rfSrc2),
    ._T_145_0(wbu__T_145_0),
    .io_in_valid_0(wbu_io_in_valid_0),
    .io_in_bits_mem_rvfi_rdata(wbu_io_in_bits_mem_rvfi_rdata),
    ._T_151_0(wbu__T_151_0),
    .io_in_bits_decode_cf_instr(wbu_io_in_bits_decode_cf_instr),
    .io_in_bits_mem_rvfi_wdata(wbu_io_in_bits_mem_rvfi_wdata),
    ._T_142_0(wbu__T_142_0),
    .io_in_bits_decode_data_src2(wbu_io_in_bits_decode_data_src2),
    .io_in_bits_mem_rvfi_rmask(wbu_io_in_bits_mem_rvfi_rmask),
    .falseWire_0(wbu_falseWire_0),
    .io_in_bits_mem_rvfi_wmask(wbu_io_in_bits_mem_rvfi_wmask)
  );
  assign io_in_0_ready = isu_io_in_0_ready; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 687:13]
  assign io_dmem_req_valid = exu_io_dmem_req_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 699:11]
  assign io_dmem_req_bits_addr = exu_io_dmem_req_bits_addr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 699:11]
  assign io_dmem_req_bits_size = exu_io_dmem_req_bits_size; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 699:11]
  assign io_dmem_req_bits_cmd = exu_io_dmem_req_bits_cmd; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 699:11]
  assign io_dmem_req_bits_wmask = exu_io_dmem_req_bits_wmask; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 699:11]
  assign io_dmem_req_bits_wdata = exu_io_dmem_req_bits_wdata; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 699:11]
  assign io_redirect_target = wbu_io__redirect_target; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 693:15]
  assign io_redirect_valid = wbu_io__redirect_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 693:15]
  assign io_in_bits_decode_data_src1 = wbu_io_in_bits_decode_data_src1;
  assign _T_2_0 = exu__T_2_0;
  assign io_in_valid = wbu_io_in_valid;
  assign io_in_bits_decode_ctrl_rfSrc1 = wbu_io_in_bits_decode_ctrl_rfSrc1;
  assign io_wb_rfDest = wbu_io_wb_rfDest;
  assign flushICache = exu_flushICache;
  assign rvfi_order = wbu_rvfi_order_0;
  assign io_in_bits_mem_rvfi_addr_real = wbu_io_in_bits_mem_rvfi_addr_real;
  assign io_in_bits_decode_ctrl_rfSrc2 = wbu_io_in_bits_decode_ctrl_rfSrc2;
  assign REG_valid = exu_REG_valid;
  assign REG_pc = exu_REG_pc;
  assign REG_isMissPredict = exu_REG_isMissPredict;
  assign REG_actualTarget = exu_REG_actualTarget;
  assign REG_actualTaken = exu_REG_actualTaken;
  assign REG_fuOpType = exu_REG_fuOpType;
  assign REG_btbType = exu_REG_btbType;
  assign REG_isRVC = exu_REG_isRVC;
  assign _T_145 = wbu__T_145_0;
  assign io_in_bits_mem_rvfi_rdata = wbu_io_in_bits_mem_rvfi_rdata;
  assign _T_151 = wbu__T_151_0;
  assign io_in_bits_decode_cf_instr = wbu_io_in_bits_decode_cf_instr;
  assign REG_0 = exu_REG_0;
  assign io_in_bits_mem_rvfi_wdata = wbu_io_in_bits_mem_rvfi_wdata;
  assign _T_142 = wbu__T_142_0;
  assign io_in_bits_decode_data_src2 = wbu_io_in_bits_decode_data_src2;
  assign intrVec = exu_intrVec;
  assign io_in_bits_mem_rvfi_rmask = wbu_io_in_bits_mem_rvfi_rmask;
  assign flushTLB = exu_flushTLB;
  assign io_in_bits_mem_rvfi_wmask = wbu_io_in_bits_mem_rvfi_wmask;
  assign isu_clock = clock;
  assign isu_reset = reset;
  assign isu_io_in_0_valid = io_in_0_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 687:13]
  assign isu_io_in_0_bits_cf_instr = io_in_0_bits_cf_instr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 687:13]
  assign isu_io_in_0_bits_cf_pc = io_in_0_bits_cf_pc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 687:13]
  assign isu_io_in_0_bits_cf_pnpc = io_in_0_bits_cf_pnpc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 687:13]
  assign isu_io_in_0_bits_cf_exceptionVec_1 = io_in_0_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 687:13]
  assign isu_io_in_0_bits_cf_exceptionVec_2 = io_in_0_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 687:13]
  assign isu_io_in_0_bits_cf_intrVec_0 = io_in_0_bits_cf_intrVec_0; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 687:13]
  assign isu_io_in_0_bits_cf_intrVec_1 = io_in_0_bits_cf_intrVec_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 687:13]
  assign isu_io_in_0_bits_cf_intrVec_2 = io_in_0_bits_cf_intrVec_2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 687:13]
  assign isu_io_in_0_bits_cf_intrVec_3 = io_in_0_bits_cf_intrVec_3; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 687:13]
  assign isu_io_in_0_bits_cf_intrVec_4 = io_in_0_bits_cf_intrVec_4; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 687:13]
  assign isu_io_in_0_bits_cf_intrVec_5 = io_in_0_bits_cf_intrVec_5; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 687:13]
  assign isu_io_in_0_bits_cf_intrVec_6 = io_in_0_bits_cf_intrVec_6; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 687:13]
  assign isu_io_in_0_bits_cf_intrVec_7 = io_in_0_bits_cf_intrVec_7; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 687:13]
  assign isu_io_in_0_bits_cf_intrVec_8 = io_in_0_bits_cf_intrVec_8; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 687:13]
  assign isu_io_in_0_bits_cf_intrVec_9 = io_in_0_bits_cf_intrVec_9; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 687:13]
  assign isu_io_in_0_bits_cf_intrVec_10 = io_in_0_bits_cf_intrVec_10; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 687:13]
  assign isu_io_in_0_bits_cf_intrVec_11 = io_in_0_bits_cf_intrVec_11; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 687:13]
  assign isu_io_in_0_bits_cf_brIdx = io_in_0_bits_cf_brIdx; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 687:13]
  assign isu_io_in_0_bits_ctrl_src1Type = io_in_0_bits_ctrl_src1Type; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 687:13]
  assign isu_io_in_0_bits_ctrl_src2Type = io_in_0_bits_ctrl_src2Type; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 687:13]
  assign isu_io_in_0_bits_ctrl_fuType = io_in_0_bits_ctrl_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 687:13]
  assign isu_io_in_0_bits_ctrl_fuOpType = io_in_0_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 687:13]
  assign isu_io_in_0_bits_ctrl_rfSrc1 = io_in_0_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 687:13]
  assign isu_io_in_0_bits_ctrl_rfSrc2 = io_in_0_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 687:13]
  assign isu_io_in_0_bits_ctrl_rfWen = io_in_0_bits_ctrl_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 687:13]
  assign isu_io_in_0_bits_ctrl_rfDest = io_in_0_bits_ctrl_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 687:13]
  assign isu_io_in_0_bits_data_imm = io_in_0_bits_data_imm; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 687:13]
  assign isu_io_out_ready = exu_io_in_ready; // @[src/main/scala/utils/Pipeline.scala 29:16]
  assign isu_io_wb_rfWen = wbu_io__wb_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 692:13]
  assign isu_io_wb_rfDest = wbu_io__wb_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 692:13]
  assign isu_io_wb_rfData = wbu_io__wb_rfData; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 692:13]
  assign isu_io_forward_valid = exu_io_forward_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 695:18]
  assign isu_io_forward_wb_rfWen = exu_io_forward_wb_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 695:18]
  assign isu_io_forward_wb_rfDest = exu_io_forward_wb_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 695:18]
  assign isu_io_forward_wb_rfData = exu_io_forward_wb_rfData; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 695:18]
  assign isu_io_forward_fuType = exu_io_forward_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 695:18]
  assign isu_io_flush = io_flush[0]; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 689:27]
  assign exu_clock = clock;
  assign exu_reset = reset;
  assign exu_io_in_valid = valid; // @[src/main/scala/utils/Pipeline.scala 31:17]
  assign exu_io_in_bits_cf_instr = exu_io_in_bits_r_cf_instr; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io_in_bits_cf_pc = exu_io_in_bits_r_cf_pc; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io_in_bits_cf_pnpc = exu_io_in_bits_r_cf_pnpc; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io_in_bits_cf_exceptionVec_1 = exu_io_in_bits_r_cf_exceptionVec_1; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io_in_bits_cf_exceptionVec_2 = exu_io_in_bits_r_cf_exceptionVec_2; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io_in_bits_cf_intrVec_0 = exu_io_in_bits_r_cf_intrVec_0; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io_in_bits_cf_intrVec_1 = exu_io_in_bits_r_cf_intrVec_1; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io_in_bits_cf_intrVec_2 = exu_io_in_bits_r_cf_intrVec_2; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io_in_bits_cf_intrVec_3 = exu_io_in_bits_r_cf_intrVec_3; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io_in_bits_cf_intrVec_4 = exu_io_in_bits_r_cf_intrVec_4; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io_in_bits_cf_intrVec_5 = exu_io_in_bits_r_cf_intrVec_5; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io_in_bits_cf_intrVec_6 = exu_io_in_bits_r_cf_intrVec_6; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io_in_bits_cf_intrVec_7 = exu_io_in_bits_r_cf_intrVec_7; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io_in_bits_cf_intrVec_8 = exu_io_in_bits_r_cf_intrVec_8; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io_in_bits_cf_intrVec_9 = exu_io_in_bits_r_cf_intrVec_9; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io_in_bits_cf_intrVec_10 = exu_io_in_bits_r_cf_intrVec_10; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io_in_bits_cf_intrVec_11 = exu_io_in_bits_r_cf_intrVec_11; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io_in_bits_cf_brIdx = exu_io_in_bits_r_cf_brIdx; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io_in_bits_ctrl_fuType = exu_io_in_bits_r_ctrl_fuType; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io_in_bits_ctrl_fuOpType = exu_io_in_bits_r_ctrl_fuOpType; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io_in_bits_ctrl_rfSrc1 = exu_io_in_bits_r_ctrl_rfSrc1; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io_in_bits_ctrl_rfSrc2 = exu_io_in_bits_r_ctrl_rfSrc2; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io_in_bits_ctrl_rfWen = exu_io_in_bits_r_ctrl_rfWen; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io_in_bits_ctrl_rfDest = exu_io_in_bits_r_ctrl_rfDest; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io_in_bits_data_src1 = exu_io_in_bits_r_data_src1; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io_in_bits_data_src2 = exu_io_in_bits_r_data_src2; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io_in_bits_data_imm = exu_io_in_bits_r_data_imm; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io_out_ready = 1'h1; // @[src/main/scala/utils/Pipeline.scala 29:16]
  assign exu_io_flush = io_flush[1]; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 690:27]
  assign exu_io_dmem_req_ready = io_dmem_req_ready; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 699:11]
  assign exu_io_dmem_resp_valid = io_dmem_resp_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 699:11]
  assign exu_io_dmem_resp_bits_rdata = io_dmem_resp_bits_rdata; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 699:11]
  assign exu_io_in_valid_0 = wbu_io_in_valid_0;
  assign exu_falseWire = wbu_falseWire_0;
  assign wbu_clock = clock;
  assign wbu_reset = reset;
  assign wbu_io__in_valid = valid_1; // @[src/main/scala/utils/Pipeline.scala 31:17]
  assign wbu_io__in_bits_decode_cf_instr = wbu_io_in_bits_r_decode_cf_instr; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_cf_pc = wbu_io_in_bits_r_decode_cf_pc; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_cf_redirect_target = wbu_io_in_bits_r_decode_cf_redirect_target; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_cf_redirect_valid = wbu_io_in_bits_r_decode_cf_redirect_valid; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_ctrl_fuType = wbu_io_in_bits_r_decode_ctrl_fuType; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_ctrl_rfSrc1 = wbu_io_in_bits_r_decode_ctrl_rfSrc1; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_ctrl_rfSrc2 = wbu_io_in_bits_r_decode_ctrl_rfSrc2; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_ctrl_rfWen = wbu_io_in_bits_r_decode_ctrl_rfWen; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_ctrl_rfDest = wbu_io_in_bits_r_decode_ctrl_rfDest; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_data_src1 = wbu_io_in_bits_r_decode_data_src1; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_data_src2 = wbu_io_in_bits_r_decode_data_src2; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_commits_0 = wbu_io_in_bits_r_commits_0; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_commits_1 = wbu_io_in_bits_r_commits_1; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_commits_2 = wbu_io_in_bits_r_commits_2; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_commits_3 = wbu_io_in_bits_r_commits_3; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_mem_rvfi_addr_real = wbu_io_in_bits_r_mem_rvfi_addr_real; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_mem_rvfi_rmask = wbu_io_in_bits_r_mem_rvfi_rmask; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_mem_rvfi_wmask = wbu_io_in_bits_r_mem_rvfi_wmask; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_mem_rvfi_rdata = wbu_io_in_bits_r_mem_rvfi_rdata; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_mem_rvfi_wdata = wbu_io_in_bits_r_mem_rvfi_wdata; // @[src/main/scala/utils/Pipeline.scala 30:16]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/Pipeline.scala 24:24]
      valid <= 1'h0; // @[src/main/scala/utils/Pipeline.scala 24:24]
    end else if (io_flush[0]) begin // @[src/main/scala/utils/Pipeline.scala 27:20]
      valid <= 1'h0; // @[src/main/scala/utils/Pipeline.scala 27:28]
    end else begin
      valid <= _GEN_1;
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_instr <= isu_io_out_bits_cf_instr; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_pc <= isu_io_out_bits_cf_pc; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_pnpc <= isu_io_out_bits_cf_pnpc; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_exceptionVec_1 <= isu_io_out_bits_cf_exceptionVec_1; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_exceptionVec_2 <= isu_io_out_bits_cf_exceptionVec_2; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_intrVec_0 <= isu_io_out_bits_cf_intrVec_0; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_intrVec_1 <= isu_io_out_bits_cf_intrVec_1; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_intrVec_2 <= isu_io_out_bits_cf_intrVec_2; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_intrVec_3 <= isu_io_out_bits_cf_intrVec_3; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_intrVec_4 <= isu_io_out_bits_cf_intrVec_4; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_intrVec_5 <= isu_io_out_bits_cf_intrVec_5; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_intrVec_6 <= isu_io_out_bits_cf_intrVec_6; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_intrVec_7 <= isu_io_out_bits_cf_intrVec_7; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_intrVec_8 <= isu_io_out_bits_cf_intrVec_8; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_intrVec_9 <= isu_io_out_bits_cf_intrVec_9; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_intrVec_10 <= isu_io_out_bits_cf_intrVec_10; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_intrVec_11 <= isu_io_out_bits_cf_intrVec_11; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_brIdx <= isu_io_out_bits_cf_brIdx; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_ctrl_fuType <= isu_io_out_bits_ctrl_fuType; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_ctrl_fuOpType <= isu_io_out_bits_ctrl_fuOpType; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_ctrl_rfSrc1 <= isu_io_out_bits_ctrl_rfSrc1; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_ctrl_rfSrc2 <= isu_io_out_bits_ctrl_rfSrc2; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_ctrl_rfWen <= isu_io_out_bits_ctrl_rfWen; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_ctrl_rfDest <= isu_io_out_bits_ctrl_rfDest; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_data_src1 <= isu_io_out_bits_data_src1; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_data_src2 <= isu_io_out_bits_data_src2; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_data_imm <= isu_io_out_bits_data_imm; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (reset) begin // @[src/main/scala/utils/Pipeline.scala 24:24]
      valid_1 <= 1'h0; // @[src/main/scala/utils/Pipeline.scala 24:24]
    end else if (io_flush[1]) begin // @[src/main/scala/utils/Pipeline.scala 27:20]
      valid_1 <= 1'h0; // @[src/main/scala/utils/Pipeline.scala 27:28]
    end else begin
      valid_1 <= _T_4;
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_decode_cf_instr <= exu_io_out_bits_decode_cf_instr; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_decode_cf_pc <= exu_io_out_bits_decode_cf_pc; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_decode_cf_redirect_target <= exu_io_out_bits_decode_cf_redirect_target; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_decode_cf_redirect_valid <= exu_io_out_bits_decode_cf_redirect_valid; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_decode_ctrl_fuType <= exu_io_out_bits_decode_ctrl_fuType; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_decode_ctrl_rfSrc1 <= exu_io_out_bits_decode_ctrl_rfSrc1; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_decode_ctrl_rfSrc2 <= exu_io_out_bits_decode_ctrl_rfSrc2; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_decode_ctrl_rfWen <= exu_io_out_bits_decode_ctrl_rfWen; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_decode_ctrl_rfDest <= exu_io_out_bits_decode_ctrl_rfDest; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_decode_data_src1 <= exu_io_out_bits_decode_data_src1; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_decode_data_src2 <= exu_io_out_bits_decode_data_src2; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_commits_0 <= exu_io_out_bits_commits_0; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_commits_1 <= exu_io_out_bits_commits_1; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_commits_2 <= exu_io_out_bits_commits_2; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_commits_3 <= exu_io_out_bits_commits_3; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_mem_rvfi_addr_real <= exu_io_out_bits_mem_rvfi_addr_real; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_mem_rvfi_rmask <= exu_io_out_bits_mem_rvfi_rmask; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_mem_rvfi_wmask <= exu_io_out_bits_mem_rvfi_wmask; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_mem_rvfi_rdata <= exu_io_out_bits_mem_rvfi_rdata; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_mem_rvfi_wdata <= exu_io_out_bits_mem_rvfi_wdata; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  valid = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  exu_io_in_bits_r_cf_instr = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  exu_io_in_bits_r_cf_pc = _RAND_2[38:0];
  _RAND_3 = {2{`RANDOM}};
  exu_io_in_bits_r_cf_pnpc = _RAND_3[38:0];
  _RAND_4 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_exceptionVec_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_exceptionVec_2 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_2 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_3 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_4 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_5 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_6 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_7 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_8 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_9 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_10 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_11 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_brIdx = _RAND_18[3:0];
  _RAND_19 = {1{`RANDOM}};
  exu_io_in_bits_r_ctrl_fuType = _RAND_19[2:0];
  _RAND_20 = {1{`RANDOM}};
  exu_io_in_bits_r_ctrl_fuOpType = _RAND_20[6:0];
  _RAND_21 = {1{`RANDOM}};
  exu_io_in_bits_r_ctrl_rfSrc1 = _RAND_21[4:0];
  _RAND_22 = {1{`RANDOM}};
  exu_io_in_bits_r_ctrl_rfSrc2 = _RAND_22[4:0];
  _RAND_23 = {1{`RANDOM}};
  exu_io_in_bits_r_ctrl_rfWen = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  exu_io_in_bits_r_ctrl_rfDest = _RAND_24[4:0];
  _RAND_25 = {2{`RANDOM}};
  exu_io_in_bits_r_data_src1 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  exu_io_in_bits_r_data_src2 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  exu_io_in_bits_r_data_imm = _RAND_27[63:0];
  _RAND_28 = {1{`RANDOM}};
  valid_1 = _RAND_28[0:0];
  _RAND_29 = {2{`RANDOM}};
  wbu_io_in_bits_r_decode_cf_instr = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  wbu_io_in_bits_r_decode_cf_pc = _RAND_30[38:0];
  _RAND_31 = {2{`RANDOM}};
  wbu_io_in_bits_r_decode_cf_redirect_target = _RAND_31[38:0];
  _RAND_32 = {1{`RANDOM}};
  wbu_io_in_bits_r_decode_cf_redirect_valid = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  wbu_io_in_bits_r_decode_ctrl_fuType = _RAND_33[2:0];
  _RAND_34 = {1{`RANDOM}};
  wbu_io_in_bits_r_decode_ctrl_rfSrc1 = _RAND_34[4:0];
  _RAND_35 = {1{`RANDOM}};
  wbu_io_in_bits_r_decode_ctrl_rfSrc2 = _RAND_35[4:0];
  _RAND_36 = {1{`RANDOM}};
  wbu_io_in_bits_r_decode_ctrl_rfWen = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  wbu_io_in_bits_r_decode_ctrl_rfDest = _RAND_37[4:0];
  _RAND_38 = {2{`RANDOM}};
  wbu_io_in_bits_r_decode_data_src1 = _RAND_38[63:0];
  _RAND_39 = {2{`RANDOM}};
  wbu_io_in_bits_r_decode_data_src2 = _RAND_39[63:0];
  _RAND_40 = {2{`RANDOM}};
  wbu_io_in_bits_r_commits_0 = _RAND_40[63:0];
  _RAND_41 = {2{`RANDOM}};
  wbu_io_in_bits_r_commits_1 = _RAND_41[63:0];
  _RAND_42 = {2{`RANDOM}};
  wbu_io_in_bits_r_commits_2 = _RAND_42[63:0];
  _RAND_43 = {2{`RANDOM}};
  wbu_io_in_bits_r_commits_3 = _RAND_43[63:0];
  _RAND_44 = {2{`RANDOM}};
  wbu_io_in_bits_r_mem_rvfi_addr_real = _RAND_44[63:0];
  _RAND_45 = {1{`RANDOM}};
  wbu_io_in_bits_r_mem_rvfi_rmask = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  wbu_io_in_bits_r_mem_rvfi_wmask = _RAND_46[7:0];
  _RAND_47 = {2{`RANDOM}};
  wbu_io_in_bits_r_mem_rvfi_rdata = _RAND_47[63:0];
  _RAND_48 = {2{`RANDOM}};
  wbu_io_in_bits_r_mem_rvfi_wdata = _RAND_48[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LockingArbiter(
  input         clock,
  input         reset,
  output        io_in_0_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input         io_in_0_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [31:0] io_in_0_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output        io_in_1_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input         io_in_1_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [31:0] io_in_1_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [2:0]  io_in_1_bits_size, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [3:0]  io_in_1_bits_cmd, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [7:0]  io_in_1_bits_wmask, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [63:0] io_in_1_bits_wdata, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input         io_out_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output        io_out_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [31:0] io_out_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [2:0]  io_out_bits_size, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [3:0]  io_out_bits_cmd, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [7:0]  io_out_bits_wmask, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [63:0] io_out_bits_wdata, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output        io_chosen // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] lockCount_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  lockIdx; // @[src/main/scala/chisel3/util/Arbiter.scala 60:22]
  wire  locked = lockCount_value != 3'h0; // @[src/main/scala/chisel3/util/Arbiter.scala 61:34]
  wire  wantsLock = io_out_bits_cmd[0] & io_out_bits_cmd[1]; // @[src/main/scala/bus/simplebus/Crossbar.scala 92:62]
  wire  _T = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [2:0] _value_T_1 = lockCount_value + 3'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  io_chosen_choice = io_in_0_valid ? 1'h0 : 1'h1; // @[src/main/scala/chisel3/util/Arbiter.scala 103:{26,35} 101:41]
  wire  _T_2 = ~io_in_0_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 45:78]
  wire  _io_in_0_ready_T_1 = locked ? ~lockIdx : 1'h1; // @[src/main/scala/chisel3/util/Arbiter.scala 71:22]
  wire  _io_in_1_ready_T_1 = locked ? lockIdx : _T_2; // @[src/main/scala/chisel3/util/Arbiter.scala 71:22]
  assign io_in_0_ready = _io_in_0_ready_T_1 & io_out_ready; // @[src/main/scala/chisel3/util/Arbiter.scala 71:56]
  assign io_in_1_ready = _io_in_1_ready_T_1 & io_out_ready; // @[src/main/scala/chisel3/util/Arbiter.scala 71:56]
  assign io_out_valid = io_chosen ? io_in_1_valid : io_in_0_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 55:{16,16}]
  assign io_out_bits_addr = io_chosen ? io_in_1_bits_addr : io_in_0_bits_addr; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_size = io_chosen ? io_in_1_bits_size : 3'h3; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_cmd = io_chosen ? io_in_1_bits_cmd : 4'h0; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_wmask = io_chosen ? io_in_1_bits_wmask : 8'h0; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_wdata = io_chosen ? io_in_1_bits_wdata : 64'h0; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_chosen = locked ? lockIdx : io_chosen_choice; // @[src/main/scala/chisel3/util/Arbiter.scala 54:13 69:{18,30}]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      lockCount_value <= 3'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (_T & wantsLock) begin // @[src/main/scala/chisel3/util/Arbiter.scala 64:36]
      lockCount_value <= _value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (_T & wantsLock) begin // @[src/main/scala/chisel3/util/Arbiter.scala 64:36]
      lockIdx <= io_chosen; // @[src/main/scala/chisel3/util/Arbiter.scala 65:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lockCount_value = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  lockIdx = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SimpleBusCrossbarNto1(
  input         clock,
  input         reset,
  output        io_in_0_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  input         io_in_0_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  input  [31:0] io_in_0_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  output        io_in_0_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  output [63:0] io_in_0_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  output        io_in_1_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  input         io_in_1_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  input  [31:0] io_in_1_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  input  [2:0]  io_in_1_req_bits_size, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  input  [3:0]  io_in_1_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  input  [7:0]  io_in_1_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  input  [63:0] io_in_1_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  output        io_in_1_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  output [3:0]  io_in_1_resp_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  output [63:0] io_in_1_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  input         io_out_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  output        io_out_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  output [31:0] io_out_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  output [2:0]  io_out_req_bits_size, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  output [3:0]  io_out_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  output [7:0]  io_out_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  output [63:0] io_out_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  output        io_out_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  input         io_out_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  input  [3:0]  io_out_resp_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  input  [63:0] io_out_resp_bits_rdata // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  inputArb_clock; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  wire  inputArb_reset; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  wire  inputArb_io_in_0_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  wire  inputArb_io_in_0_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  wire [31:0] inputArb_io_in_0_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  wire  inputArb_io_in_1_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  wire  inputArb_io_in_1_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  wire [31:0] inputArb_io_in_1_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  wire [2:0] inputArb_io_in_1_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  wire [3:0] inputArb_io_in_1_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  wire [7:0] inputArb_io_in_1_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  wire [63:0] inputArb_io_in_1_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  wire  inputArb_io_out_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  wire  inputArb_io_out_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  wire [31:0] inputArb_io_out_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  wire [2:0] inputArb_io_out_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  wire [3:0] inputArb_io_out_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  wire [7:0] inputArb_io_out_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  wire [63:0] inputArb_io_out_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  wire  inputArb_io_chosen; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  reg [1:0] state; // @[src/main/scala/bus/simplebus/Crossbar.scala 90:22]
  reg  inflightSrc; // @[src/main/scala/bus/simplebus/Crossbar.scala 97:28]
  wire  _io_out_req_valid_T = state == 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:47]
  wire  _T_1 = inputArb_io_out_ready & inputArb_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _T_6 = ~inputArb_io_out_bits_cmd[0] & ~inputArb_io_out_bits_cmd[3]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:26]
  wire  _T_7 = inputArb_io_out_bits_cmd == 4'h7; // @[src/main/scala/bus/simplebus/SimpleBus.scala 78:27]
  wire  _T_8 = inputArb_io_out_bits_cmd == 4'h1; // @[src/main/scala/bus/simplebus/SimpleBus.scala 77:29]
  wire [1:0] _GEN_4 = _T_7 | _T_8 ? 2'h2 : state; // @[src/main/scala/bus/simplebus/Crossbar.scala 116:{80,88} 90:22]
  wire  _T_11 = io_out_resp_ready & io_out_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _T_12 = io_out_resp_bits_cmd == 4'h6; // @[src/main/scala/bus/simplebus/SimpleBus.scala 91:26]
  wire [1:0] _GEN_9 = _T_11 ? 2'h0 : state; // @[src/main/scala/bus/simplebus/Crossbar.scala 120:{48,56} 90:22]
  LockingArbiter inputArb ( // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
    .clock(inputArb_clock),
    .reset(inputArb_reset),
    .io_in_0_ready(inputArb_io_in_0_ready),
    .io_in_0_valid(inputArb_io_in_0_valid),
    .io_in_0_bits_addr(inputArb_io_in_0_bits_addr),
    .io_in_1_ready(inputArb_io_in_1_ready),
    .io_in_1_valid(inputArb_io_in_1_valid),
    .io_in_1_bits_addr(inputArb_io_in_1_bits_addr),
    .io_in_1_bits_size(inputArb_io_in_1_bits_size),
    .io_in_1_bits_cmd(inputArb_io_in_1_bits_cmd),
    .io_in_1_bits_wmask(inputArb_io_in_1_bits_wmask),
    .io_in_1_bits_wdata(inputArb_io_in_1_bits_wdata),
    .io_out_ready(inputArb_io_out_ready),
    .io_out_valid(inputArb_io_out_valid),
    .io_out_bits_addr(inputArb_io_out_bits_addr),
    .io_out_bits_size(inputArb_io_out_bits_size),
    .io_out_bits_cmd(inputArb_io_out_bits_cmd),
    .io_out_bits_wmask(inputArb_io_out_bits_wmask),
    .io_out_bits_wdata(inputArb_io_out_bits_wdata),
    .io_chosen(inputArb_io_chosen)
  );
  assign io_in_0_req_ready = inputArb_io_in_0_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 94:68]
  assign io_in_0_resp_valid = ~inflightSrc & io_out_resp_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 107:{13,13} 105:26]
  assign io_in_0_resp_bits_rdata = io_out_resp_bits_rdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 104:25]
  assign io_in_1_req_ready = inputArb_io_in_1_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 94:68]
  assign io_in_1_resp_valid = inflightSrc & io_out_resp_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 107:{13,13} 105:26]
  assign io_in_1_resp_bits_cmd = io_out_resp_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 104:25]
  assign io_in_1_resp_bits_rdata = io_out_resp_bits_rdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 104:25]
  assign io_out_req_valid = inputArb_io_out_valid & state == 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:37]
  assign io_out_req_bits_addr = inputArb_io_out_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 99:19]
  assign io_out_req_bits_size = inputArb_io_out_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 99:19]
  assign io_out_req_bits_cmd = inputArb_io_out_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 99:19]
  assign io_out_req_bits_wmask = inputArb_io_out_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 99:19]
  assign io_out_req_bits_wdata = inputArb_io_out_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 99:19]
  assign io_out_resp_ready = 1'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 108:{13,13}]
  assign inputArb_clock = clock;
  assign inputArb_reset = reset;
  assign inputArb_io_in_0_valid = io_in_0_req_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 94:68]
  assign inputArb_io_in_0_bits_addr = io_in_0_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 94:68]
  assign inputArb_io_in_1_valid = io_in_1_req_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 94:68]
  assign inputArb_io_in_1_bits_addr = io_in_1_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 94:68]
  assign inputArb_io_in_1_bits_size = io_in_1_req_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 94:68]
  assign inputArb_io_in_1_bits_cmd = io_in_1_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 94:68]
  assign inputArb_io_in_1_bits_wmask = io_in_1_req_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 94:68]
  assign inputArb_io_in_1_bits_wdata = io_in_1_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 94:68]
  assign inputArb_io_out_ready = io_out_req_ready & _io_out_req_valid_T; // @[src/main/scala/bus/simplebus/Crossbar.scala 102:37]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 90:22]
      state <= 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 90:22]
    end else if (2'h0 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 111:18]
      if (_T_1) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:27]
        if (_T_6) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 115:38]
          state <= 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 115:46]
        end else begin
          state <= _GEN_4;
        end
      end
    end else if (2'h1 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 111:18]
      if (_T_11 & _T_12) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 119:80]
        state <= 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 119:88]
      end
    end else if (2'h2 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 111:18]
      state <= _GEN_9;
    end
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 97:28]
      inflightSrc <= 1'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 97:28]
    end else if (2'h0 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 111:18]
      if (_T_1) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:27]
        inflightSrc <= inputArb_io_chosen; // @[src/main/scala/bus/simplebus/Crossbar.scala 114:21]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  inflightSrc = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LockingArbiter_1(
  input         clock,
  input         reset,
  output        io_in_0_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input         io_in_0_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [31:0] io_in_0_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [2:0]  io_in_0_bits_size, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [3:0]  io_in_0_bits_cmd, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [7:0]  io_in_0_bits_wmask, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [63:0] io_in_0_bits_wdata, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output        io_in_3_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input         io_in_3_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [31:0] io_in_3_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [2:0]  io_in_3_bits_size, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [3:0]  io_in_3_bits_cmd, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [7:0]  io_in_3_bits_wmask, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [63:0] io_in_3_bits_wdata, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input         io_out_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output        io_out_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [31:0] io_out_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [2:0]  io_out_bits_size, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [3:0]  io_out_bits_cmd, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [7:0]  io_out_bits_wmask, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [63:0] io_out_bits_wdata, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [1:0]  io_chosen // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  _GEN_1 = 2'h1 == io_chosen ? 1'h0 : io_in_0_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 55:{16,16}]
  wire  _GEN_2 = 2'h2 == io_chosen ? 1'h0 : _GEN_1; // @[src/main/scala/chisel3/util/Arbiter.scala 55:{16,16}]
  wire [31:0] _GEN_5 = 2'h1 == io_chosen ? 32'h0 : io_in_0_bits_addr; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire [31:0] _GEN_6 = 2'h2 == io_chosen ? 32'h0 : _GEN_5; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire [2:0] _GEN_9 = 2'h1 == io_chosen ? 3'h0 : io_in_0_bits_size; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire [2:0] _GEN_10 = 2'h2 == io_chosen ? 3'h0 : _GEN_9; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire [3:0] _GEN_13 = 2'h1 == io_chosen ? 4'h0 : io_in_0_bits_cmd; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire [3:0] _GEN_14 = 2'h2 == io_chosen ? 4'h0 : _GEN_13; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire [7:0] _GEN_17 = 2'h1 == io_chosen ? 8'h0 : io_in_0_bits_wmask; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire [7:0] _GEN_18 = 2'h2 == io_chosen ? 8'h0 : _GEN_17; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire [63:0] _GEN_21 = 2'h1 == io_chosen ? 64'h0 : io_in_0_bits_wdata; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire [63:0] _GEN_22 = 2'h2 == io_chosen ? 64'h0 : _GEN_21; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  reg [2:0] lockCount_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg [1:0] lockIdx; // @[src/main/scala/chisel3/util/Arbiter.scala 60:22]
  wire  locked = lockCount_value != 3'h0; // @[src/main/scala/chisel3/util/Arbiter.scala 61:34]
  wire  wantsLock = io_out_bits_cmd[0] & io_out_bits_cmd[1]; // @[src/main/scala/bus/simplebus/Crossbar.scala 92:62]
  wire  _T = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [2:0] _value_T_1 = lockCount_value + 3'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire [1:0] io_chosen_choice = io_in_0_valid ? 2'h0 : 2'h3; // @[src/main/scala/chisel3/util/Arbiter.scala 103:{26,35}]
  wire  _T_4 = ~io_in_0_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 45:78]
  wire  _io_in_0_ready_T_1 = locked ? lockIdx == 2'h0 : 1'h1; // @[src/main/scala/chisel3/util/Arbiter.scala 71:22]
  wire  _io_in_3_ready_T_1 = locked ? lockIdx == 2'h3 : _T_4; // @[src/main/scala/chisel3/util/Arbiter.scala 71:22]
  assign io_in_0_ready = _io_in_0_ready_T_1 & io_out_ready; // @[src/main/scala/chisel3/util/Arbiter.scala 71:56]
  assign io_in_3_ready = _io_in_3_ready_T_1 & io_out_ready; // @[src/main/scala/chisel3/util/Arbiter.scala 71:56]
  assign io_out_valid = 2'h3 == io_chosen ? io_in_3_valid : _GEN_2; // @[src/main/scala/chisel3/util/Arbiter.scala 55:{16,16}]
  assign io_out_bits_addr = 2'h3 == io_chosen ? io_in_3_bits_addr : _GEN_6; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_size = 2'h3 == io_chosen ? io_in_3_bits_size : _GEN_10; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_cmd = 2'h3 == io_chosen ? io_in_3_bits_cmd : _GEN_14; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_wmask = 2'h3 == io_chosen ? io_in_3_bits_wmask : _GEN_18; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_wdata = 2'h3 == io_chosen ? io_in_3_bits_wdata : _GEN_22; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_chosen = locked ? lockIdx : io_chosen_choice; // @[src/main/scala/chisel3/util/Arbiter.scala 54:13 69:{18,30}]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      lockCount_value <= 3'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (_T & wantsLock) begin // @[src/main/scala/chisel3/util/Arbiter.scala 64:36]
      lockCount_value <= _value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (_T & wantsLock) begin // @[src/main/scala/chisel3/util/Arbiter.scala 64:36]
      lockIdx <= io_chosen; // @[src/main/scala/chisel3/util/Arbiter.scala 65:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lockCount_value = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  lockIdx = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SimpleBusCrossbarNto1_1(
  input         clock,
  input         reset,
  output        io_in_0_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  input         io_in_0_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  input  [31:0] io_in_0_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  input  [2:0]  io_in_0_req_bits_size, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  input  [3:0]  io_in_0_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  input  [7:0]  io_in_0_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  input  [63:0] io_in_0_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  output        io_in_0_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  output [63:0] io_in_0_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  output        io_in_3_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  input         io_in_3_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  input  [31:0] io_in_3_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  input  [2:0]  io_in_3_req_bits_size, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  input  [3:0]  io_in_3_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  input  [7:0]  io_in_3_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  input  [63:0] io_in_3_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  input         io_in_3_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  output        io_in_3_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  output [3:0]  io_in_3_resp_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  output [63:0] io_in_3_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  input         io_out_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  output        io_out_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  output [31:0] io_out_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  output [2:0]  io_out_req_bits_size, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  output [3:0]  io_out_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  output [7:0]  io_out_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  output [63:0] io_out_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  output        io_out_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  input         io_out_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  input  [3:0]  io_out_resp_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
  input  [63:0] io_out_resp_bits_rdata // @[src/main/scala/bus/simplebus/Crossbar.scala 84:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  inputArb_clock; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  wire  inputArb_reset; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  wire  inputArb_io_in_0_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  wire  inputArb_io_in_0_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  wire [31:0] inputArb_io_in_0_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  wire [2:0] inputArb_io_in_0_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  wire [3:0] inputArb_io_in_0_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  wire [7:0] inputArb_io_in_0_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  wire [63:0] inputArb_io_in_0_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  wire  inputArb_io_in_3_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  wire  inputArb_io_in_3_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  wire [31:0] inputArb_io_in_3_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  wire [2:0] inputArb_io_in_3_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  wire [3:0] inputArb_io_in_3_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  wire [7:0] inputArb_io_in_3_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  wire [63:0] inputArb_io_in_3_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  wire  inputArb_io_out_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  wire  inputArb_io_out_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  wire [31:0] inputArb_io_out_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  wire [2:0] inputArb_io_out_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  wire [3:0] inputArb_io_out_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  wire [7:0] inputArb_io_out_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  wire [63:0] inputArb_io_out_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  wire [1:0] inputArb_io_chosen; // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
  reg [1:0] state; // @[src/main/scala/bus/simplebus/Crossbar.scala 90:22]
  reg [1:0] inflightSrc; // @[src/main/scala/bus/simplebus/Crossbar.scala 97:28]
  wire  _io_out_req_valid_T = state == 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:47]
  wire  _GEN_5 = 2'h1 == inflightSrc ? 1'h0 : 1'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 108:{13,13}]
  wire  _GEN_6 = 2'h2 == inflightSrc ? 1'h0 : _GEN_5; // @[src/main/scala/bus/simplebus/Crossbar.scala 108:{13,13}]
  wire  _T_1 = inputArb_io_out_ready & inputArb_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _T_6 = ~inputArb_io_out_bits_cmd[0] & ~inputArb_io_out_bits_cmd[3]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:26]
  wire  _T_7 = inputArb_io_out_bits_cmd == 4'h7; // @[src/main/scala/bus/simplebus/SimpleBus.scala 78:27]
  wire  _T_8 = inputArb_io_out_bits_cmd == 4'h1; // @[src/main/scala/bus/simplebus/SimpleBus.scala 77:29]
  wire [1:0] _GEN_8 = _T_7 | _T_8 ? 2'h2 : state; // @[src/main/scala/bus/simplebus/Crossbar.scala 116:{80,88} 90:22]
  wire  _T_11 = io_out_resp_ready & io_out_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _T_12 = io_out_resp_bits_cmd == 4'h6; // @[src/main/scala/bus/simplebus/SimpleBus.scala 91:26]
  wire [1:0] _GEN_13 = _T_11 ? 2'h0 : state; // @[src/main/scala/bus/simplebus/Crossbar.scala 120:{48,56} 90:22]
  LockingArbiter_1 inputArb ( // @[src/main/scala/bus/simplebus/Crossbar.scala 93:24]
    .clock(inputArb_clock),
    .reset(inputArb_reset),
    .io_in_0_ready(inputArb_io_in_0_ready),
    .io_in_0_valid(inputArb_io_in_0_valid),
    .io_in_0_bits_addr(inputArb_io_in_0_bits_addr),
    .io_in_0_bits_size(inputArb_io_in_0_bits_size),
    .io_in_0_bits_cmd(inputArb_io_in_0_bits_cmd),
    .io_in_0_bits_wmask(inputArb_io_in_0_bits_wmask),
    .io_in_0_bits_wdata(inputArb_io_in_0_bits_wdata),
    .io_in_3_ready(inputArb_io_in_3_ready),
    .io_in_3_valid(inputArb_io_in_3_valid),
    .io_in_3_bits_addr(inputArb_io_in_3_bits_addr),
    .io_in_3_bits_size(inputArb_io_in_3_bits_size),
    .io_in_3_bits_cmd(inputArb_io_in_3_bits_cmd),
    .io_in_3_bits_wmask(inputArb_io_in_3_bits_wmask),
    .io_in_3_bits_wdata(inputArb_io_in_3_bits_wdata),
    .io_out_ready(inputArb_io_out_ready),
    .io_out_valid(inputArb_io_out_valid),
    .io_out_bits_addr(inputArb_io_out_bits_addr),
    .io_out_bits_size(inputArb_io_out_bits_size),
    .io_out_bits_cmd(inputArb_io_out_bits_cmd),
    .io_out_bits_wmask(inputArb_io_out_bits_wmask),
    .io_out_bits_wdata(inputArb_io_out_bits_wdata),
    .io_chosen(inputArb_io_chosen)
  );
  assign io_in_0_req_ready = inputArb_io_in_0_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 94:68]
  assign io_in_0_resp_valid = 2'h0 == inflightSrc & io_out_resp_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 107:{13,13} 105:26]
  assign io_in_0_resp_bits_rdata = io_out_resp_bits_rdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 104:25]
  assign io_in_3_req_ready = inputArb_io_in_3_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 94:68]
  assign io_in_3_resp_valid = 2'h3 == inflightSrc & io_out_resp_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 107:{13,13} 105:26]
  assign io_in_3_resp_bits_cmd = io_out_resp_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 104:25]
  assign io_in_3_resp_bits_rdata = io_out_resp_bits_rdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 104:25]
  assign io_out_req_valid = inputArb_io_out_valid & state == 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:37]
  assign io_out_req_bits_addr = inputArb_io_out_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 99:19]
  assign io_out_req_bits_size = inputArb_io_out_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 99:19]
  assign io_out_req_bits_cmd = inputArb_io_out_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 99:19]
  assign io_out_req_bits_wmask = inputArb_io_out_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 99:19]
  assign io_out_req_bits_wdata = inputArb_io_out_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 99:19]
  assign io_out_resp_ready = 2'h3 == inflightSrc ? io_in_3_resp_ready : _GEN_6; // @[src/main/scala/bus/simplebus/Crossbar.scala 108:{13,13}]
  assign inputArb_clock = clock;
  assign inputArb_reset = reset;
  assign inputArb_io_in_0_valid = io_in_0_req_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 94:68]
  assign inputArb_io_in_0_bits_addr = io_in_0_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 94:68]
  assign inputArb_io_in_0_bits_size = io_in_0_req_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 94:68]
  assign inputArb_io_in_0_bits_cmd = io_in_0_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 94:68]
  assign inputArb_io_in_0_bits_wmask = io_in_0_req_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 94:68]
  assign inputArb_io_in_0_bits_wdata = io_in_0_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 94:68]
  assign inputArb_io_in_3_valid = io_in_3_req_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 94:68]
  assign inputArb_io_in_3_bits_addr = io_in_3_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 94:68]
  assign inputArb_io_in_3_bits_size = io_in_3_req_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 94:68]
  assign inputArb_io_in_3_bits_cmd = io_in_3_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 94:68]
  assign inputArb_io_in_3_bits_wmask = io_in_3_req_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 94:68]
  assign inputArb_io_in_3_bits_wdata = io_in_3_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 94:68]
  assign inputArb_io_out_ready = io_out_req_ready & _io_out_req_valid_T; // @[src/main/scala/bus/simplebus/Crossbar.scala 102:37]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 90:22]
      state <= 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 90:22]
    end else if (2'h0 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 111:18]
      if (_T_1) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:27]
        if (_T_6) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 115:38]
          state <= 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 115:46]
        end else begin
          state <= _GEN_8;
        end
      end
    end else if (2'h1 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 111:18]
      if (_T_11 & _T_12) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 119:80]
        state <= 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 119:88]
      end
    end else if (2'h2 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 111:18]
      state <= _GEN_13;
    end
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 97:28]
      inflightSrc <= 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 97:28]
    end else if (2'h0 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 111:18]
      if (_T_1) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:27]
        inflightSrc <= inputArb_io_chosen; // @[src/main/scala/bus/simplebus/Crossbar.scala 114:21]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  inflightSrc = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module EmbeddedTLB_fake(
  output        io_in_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 39:14]
  input         io_in_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 39:14]
  input  [38:0] io_in_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 39:14]
  input  [86:0] io_in_req_bits_user, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 39:14]
  input         io_in_resp_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 39:14]
  output        io_in_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 39:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 39:14]
  output [86:0] io_in_resp_bits_user, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 39:14]
  input         io_out_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 39:14]
  output        io_out_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 39:14]
  output [31:0] io_out_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 39:14]
  output [86:0] io_out_req_bits_user, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 39:14]
  output        io_out_resp_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 39:14]
  input         io_out_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 39:14]
  input  [63:0] io_out_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 39:14]
  input  [86:0] io_out_resp_bits_user // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 39:14]
);
  assign io_in_req_ready = io_out_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 425:10]
  assign io_in_resp_valid = io_out_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 425:10]
  assign io_in_resp_bits_rdata = io_out_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 425:10]
  assign io_in_resp_bits_user = io_out_resp_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 425:10]
  assign io_out_req_valid = io_in_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 425:10]
  assign io_out_req_bits_addr = io_in_req_bits_addr[31:0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 425:10]
  assign io_out_req_bits_user = io_in_req_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 425:10]
  assign io_out_resp_ready = io_in_resp_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 425:10]
endmodule
module Cache_fake(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_in_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [86:0] io_in_req_bits_user, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_in_resp_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output        io_in_resp_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [86:0] io_in_resp_bits_user, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [1:0]  io_flush, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_out_mem_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output        io_out_mem_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [31:0] io_out_mem_req_bits_addr, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output        io_out_mem_resp_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_out_mem_resp_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [63:0] io_out_mem_resp_bits_rdata, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_mmio_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output        io_mmio_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [31:0] io_mmio_req_bits_addr, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output        io_mmio_resp_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_mmio_resp_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [63:0] io_mmio_resp_bits_rdata // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [95:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[src/main/scala/nutcore/mem/Cache.scala 558:22]
  wire [31:0] _ismmio_T = io_in_req_bits_addr ^ 32'h30000000; // @[src/main/scala/nutcore/NutCore.scala 103:11]
  wire  _ismmio_T_2 = _ismmio_T[31:28] == 4'h0; // @[src/main/scala/nutcore/NutCore.scala 103:44]
  wire [31:0] _ismmio_T_3 = io_in_req_bits_addr ^ 32'h40000000; // @[src/main/scala/nutcore/NutCore.scala 103:11]
  wire  _ismmio_T_5 = _ismmio_T_3[31:30] == 2'h0; // @[src/main/scala/nutcore/NutCore.scala 103:44]
  wire  ismmio = _ismmio_T_2 | _ismmio_T_5; // @[src/main/scala/nutcore/NutCore.scala 104:15]
  wire  _ismmioRec_T = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  ismmioRec; // @[src/main/scala/nutcore/mem/Cache.scala 561:28]
  reg  needFlush; // @[src/main/scala/nutcore/mem/Cache.scala 566:26]
  wire  _GEN_1 = io_flush[0] & state != 3'h0 | needFlush; // @[src/main/scala/nutcore/mem/Cache.scala 566:26 567:{44,56}]
  wire  _alreadyOutFire_T = io_in_resp_ready & io_in_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  alreadyOutFire; // @[src/main/scala/nutcore/mem/Cache.scala 570:33]
  wire  _GEN_3 = _alreadyOutFire_T | alreadyOutFire; // @[src/main/scala/nutcore/mem/Cache.scala 570:{33,33,33}]
  wire  _T_11 = io_out_mem_req_ready & io_out_mem_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _T_13 = io_out_mem_resp_ready & io_out_mem_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [2:0] _GEN_6 = _T_13 ? 3'h5 : state; // @[src/main/scala/nutcore/mem/Cache.scala 558:22 581:{35,43}]
  wire  _T_15 = io_mmio_req_ready & io_mmio_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [2:0] _GEN_7 = _T_15 ? 3'h4 : state; // @[src/main/scala/nutcore/mem/Cache.scala 558:22 584:{31,39}]
  wire  _T_17 = io_mmio_resp_ready & io_mmio_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [2:0] _GEN_8 = _T_17 | alreadyOutFire ? 3'h5 : state; // @[src/main/scala/nutcore/mem/Cache.scala 558:22 587:{50,58}]
  wire [2:0] _GEN_9 = _alreadyOutFire_T | needFlush | alreadyOutFire ? 3'h0 : state; // @[src/main/scala/nutcore/mem/Cache.scala 558:22 590:{61,69}]
  wire [2:0] _GEN_10 = 3'h5 == state ? _GEN_9 : state; // @[src/main/scala/nutcore/mem/Cache.scala 572:18 558:22]
  wire [2:0] _GEN_11 = 3'h4 == state ? _GEN_8 : _GEN_10; // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
  wire [2:0] _GEN_12 = 3'h3 == state ? _GEN_7 : _GEN_11; // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
  reg [31:0] reqaddr; // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
  reg [63:0] mmiordata; // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
  reg [63:0] memrdata; // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
  reg [86:0] memuser; // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
  assign io_in_req_ready = state == 3'h0; // @[src/main/scala/nutcore/mem/Cache.scala 600:29]
  assign io_in_resp_valid = state == 3'h5 & ~needFlush; // @[src/main/scala/nutcore/mem/Cache.scala 601:47]
  assign io_in_resp_bits_rdata = ismmioRec ? mmiordata : memrdata; // @[src/main/scala/nutcore/mem/Cache.scala 608:31]
  assign io_in_resp_bits_user = memuser; // @[src/main/scala/nutcore/mem/Cache.scala 612:93]
  assign io_out_mem_req_valid = state == 3'h1; // @[src/main/scala/nutcore/mem/Cache.scala 617:34]
  assign io_out_mem_req_bits_addr = reqaddr; // @[src/main/scala/bus/simplebus/SimpleBus.scala 64:15]
  assign io_out_mem_resp_ready = 1'h1; // @[src/main/scala/nutcore/mem/Cache.scala 618:25]
  assign io_mmio_req_valid = state == 3'h3; // @[src/main/scala/nutcore/mem/Cache.scala 623:31]
  assign io_mmio_req_bits_addr = reqaddr; // @[src/main/scala/bus/simplebus/SimpleBus.scala 64:15]
  assign io_mmio_resp_ready = 1'h1; // @[src/main/scala/nutcore/mem/Cache.scala 624:22]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/mem/Cache.scala 558:22]
      state <= 3'h0; // @[src/main/scala/nutcore/mem/Cache.scala 558:22]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
      if (_ismmioRec_T & ~io_flush[0]) begin // @[src/main/scala/nutcore/mem/Cache.scala 575:45]
        if (ismmio) begin // @[src/main/scala/nutcore/mem/Cache.scala 575:59]
          state <= 3'h3;
        end else begin
          state <= 3'h1;
        end
      end
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
      if (_T_11) begin // @[src/main/scala/nutcore/mem/Cache.scala 578:34]
        state <= 3'h2; // @[src/main/scala/nutcore/mem/Cache.scala 578:42]
      end
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
      state <= _GEN_6;
    end else begin
      state <= _GEN_12;
    end
    if (_ismmioRec_T) begin // @[src/main/scala/nutcore/mem/Cache.scala 561:28]
      ismmioRec <= ismmio; // @[src/main/scala/nutcore/mem/Cache.scala 561:28]
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/Cache.scala 566:26]
      needFlush <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 566:26]
    end else if (state == 3'h0 & needFlush) begin // @[src/main/scala/nutcore/mem/Cache.scala 568:40]
      needFlush <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 568:52]
    end else begin
      needFlush <= _GEN_1;
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/Cache.scala 570:33]
      alreadyOutFire <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 570:33]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
      alreadyOutFire <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 574:22]
    end else begin
      alreadyOutFire <= _GEN_3;
    end
    if (_ismmioRec_T) begin // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
      reqaddr <= io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    if (_T_17) begin // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
      mmiordata <= io_mmio_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    if (_T_13) begin // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
      memrdata <= io_out_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    if (_ismmioRec_T) begin // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
      memuser <= io_in_req_bits_user; // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  ismmioRec = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  needFlush = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  alreadyOutFire = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  reqaddr = _RAND_4[31:0];
  _RAND_5 = {2{`RANDOM}};
  mmiordata = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  memrdata = _RAND_6[63:0];
  _RAND_7 = {3{`RANDOM}};
  memuser = _RAND_7[86:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module EmbeddedTLB_fake_1(
  output        io_in_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 39:14]
  input         io_in_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 39:14]
  input  [38:0] io_in_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 39:14]
  input  [2:0]  io_in_req_bits_size, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 39:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 39:14]
  input  [7:0]  io_in_req_bits_wmask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 39:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 39:14]
  output        io_in_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 39:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 39:14]
  input         io_out_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 39:14]
  output        io_out_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 39:14]
  output [31:0] io_out_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 39:14]
  output [2:0]  io_out_req_bits_size, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 39:14]
  output [3:0]  io_out_req_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 39:14]
  output [7:0]  io_out_req_bits_wmask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 39:14]
  output [63:0] io_out_req_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 39:14]
  input         io_out_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 39:14]
  input  [63:0] io_out_resp_bits_rdata // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 39:14]
);
  assign io_in_req_ready = io_out_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 425:10]
  assign io_in_resp_valid = io_out_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 425:10]
  assign io_in_resp_bits_rdata = io_out_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 425:10]
  assign io_out_req_valid = io_in_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 425:10]
  assign io_out_req_bits_addr = io_in_req_bits_addr[31:0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 425:10]
  assign io_out_req_bits_size = io_in_req_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 425:10]
  assign io_out_req_bits_cmd = io_in_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 425:10]
  assign io_out_req_bits_wmask = io_in_req_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 425:10]
  assign io_out_req_bits_wdata = io_in_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 425:10]
endmodule
module Cache_fake_1(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_in_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [2:0]  io_in_req_bits_size, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [7:0]  io_in_req_bits_wmask, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_in_resp_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output        io_in_resp_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [3:0]  io_in_resp_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_out_mem_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output        io_out_mem_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [31:0] io_out_mem_req_bits_addr, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [2:0]  io_out_mem_req_bits_size, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [3:0]  io_out_mem_req_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [7:0]  io_out_mem_req_bits_wmask, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [63:0] io_out_mem_req_bits_wdata, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output        io_out_mem_resp_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_out_mem_resp_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [3:0]  io_out_mem_resp_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [63:0] io_out_mem_resp_bits_rdata, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_mmio_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output        io_mmio_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [31:0] io_mmio_req_bits_addr, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [2:0]  io_mmio_req_bits_size, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [3:0]  io_mmio_req_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [7:0]  io_mmio_req_bits_wmask, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [63:0] io_mmio_req_bits_wdata, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output        io_mmio_resp_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_mmio_resp_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [3:0]  io_mmio_resp_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [63:0] io_mmio_resp_bits_rdata // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[src/main/scala/nutcore/mem/Cache.scala 558:22]
  wire [31:0] _ismmio_T = io_in_req_bits_addr ^ 32'h30000000; // @[src/main/scala/nutcore/NutCore.scala 103:11]
  wire  _ismmio_T_2 = _ismmio_T[31:28] == 4'h0; // @[src/main/scala/nutcore/NutCore.scala 103:44]
  wire [31:0] _ismmio_T_3 = io_in_req_bits_addr ^ 32'h40000000; // @[src/main/scala/nutcore/NutCore.scala 103:11]
  wire  _ismmio_T_5 = _ismmio_T_3[31:30] == 2'h0; // @[src/main/scala/nutcore/NutCore.scala 103:44]
  wire  ismmio = _ismmio_T_2 | _ismmio_T_5; // @[src/main/scala/nutcore/NutCore.scala 104:15]
  wire  _ismmioRec_T = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  ismmioRec; // @[src/main/scala/nutcore/mem/Cache.scala 561:28]
  wire  _alreadyOutFire_T = io_in_resp_ready & io_in_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  reg  alreadyOutFire; // @[src/main/scala/nutcore/mem/Cache.scala 570:33]
  wire  _GEN_3 = _alreadyOutFire_T | alreadyOutFire; // @[src/main/scala/nutcore/mem/Cache.scala 570:{33,33,33}]
  wire  _T_11 = io_out_mem_req_ready & io_out_mem_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire  _T_13 = io_out_mem_resp_ready & io_out_mem_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [2:0] _GEN_6 = _T_13 ? 3'h5 : state; // @[src/main/scala/nutcore/mem/Cache.scala 558:22 581:{35,43}]
  wire  _T_15 = io_mmio_req_ready & io_mmio_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [2:0] _GEN_7 = _T_15 ? 3'h4 : state; // @[src/main/scala/nutcore/mem/Cache.scala 558:22 584:{31,39}]
  wire  _T_17 = io_mmio_resp_ready & io_mmio_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [2:0] _GEN_8 = _T_17 | alreadyOutFire ? 3'h5 : state; // @[src/main/scala/nutcore/mem/Cache.scala 558:22 587:{50,58}]
  wire [2:0] _GEN_9 = _GEN_3 ? 3'h0 : state; // @[src/main/scala/nutcore/mem/Cache.scala 558:22 590:{61,69}]
  wire [2:0] _GEN_10 = 3'h5 == state ? _GEN_9 : state; // @[src/main/scala/nutcore/mem/Cache.scala 572:18 558:22]
  wire [2:0] _GEN_11 = 3'h4 == state ? _GEN_8 : _GEN_10; // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
  wire [2:0] _GEN_12 = 3'h3 == state ? _GEN_7 : _GEN_11; // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
  reg [31:0] reqaddr; // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
  reg [3:0] cmd; // @[src/main/scala/nutcore/mem/Cache.scala 595:22]
  reg [2:0] size; // @[src/main/scala/nutcore/mem/Cache.scala 596:23]
  reg [63:0] wdata; // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
  reg [7:0] wmask; // @[src/main/scala/nutcore/mem/Cache.scala 598:24]
  reg [63:0] mmiordata; // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
  reg [3:0] mmiocmd; // @[src/main/scala/nutcore/mem/Cache.scala 604:26]
  reg [63:0] memrdata; // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
  reg [3:0] memcmd; // @[src/main/scala/nutcore/mem/Cache.scala 606:25]
  assign io_in_req_ready = state == 3'h0; // @[src/main/scala/nutcore/mem/Cache.scala 600:29]
  assign io_in_resp_valid = state == 3'h5; // @[src/main/scala/nutcore/mem/Cache.scala 601:30]
  assign io_in_resp_bits_cmd = ismmioRec ? mmiocmd : memcmd; // @[src/main/scala/nutcore/mem/Cache.scala 609:29]
  assign io_in_resp_bits_rdata = ismmioRec ? mmiordata : memrdata; // @[src/main/scala/nutcore/mem/Cache.scala 608:31]
  assign io_out_mem_req_valid = state == 3'h1; // @[src/main/scala/nutcore/mem/Cache.scala 617:34]
  assign io_out_mem_req_bits_addr = reqaddr; // @[src/main/scala/bus/simplebus/SimpleBus.scala 64:15]
  assign io_out_mem_req_bits_size = size; // @[src/main/scala/bus/simplebus/SimpleBus.scala 66:15]
  assign io_out_mem_req_bits_cmd = cmd; // @[src/main/scala/bus/simplebus/SimpleBus.scala 65:14]
  assign io_out_mem_req_bits_wmask = wmask; // @[src/main/scala/bus/simplebus/SimpleBus.scala 68:16]
  assign io_out_mem_req_bits_wdata = wdata; // @[src/main/scala/bus/simplebus/SimpleBus.scala 67:16]
  assign io_out_mem_resp_ready = 1'h1; // @[src/main/scala/nutcore/mem/Cache.scala 618:25]
  assign io_mmio_req_valid = state == 3'h3; // @[src/main/scala/nutcore/mem/Cache.scala 623:31]
  assign io_mmio_req_bits_addr = reqaddr; // @[src/main/scala/bus/simplebus/SimpleBus.scala 64:15]
  assign io_mmio_req_bits_size = size; // @[src/main/scala/bus/simplebus/SimpleBus.scala 66:15]
  assign io_mmio_req_bits_cmd = cmd; // @[src/main/scala/bus/simplebus/SimpleBus.scala 65:14]
  assign io_mmio_req_bits_wmask = wmask; // @[src/main/scala/bus/simplebus/SimpleBus.scala 68:16]
  assign io_mmio_req_bits_wdata = wdata; // @[src/main/scala/bus/simplebus/SimpleBus.scala 67:16]
  assign io_mmio_resp_ready = 1'h1; // @[src/main/scala/nutcore/mem/Cache.scala 624:22]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/mem/Cache.scala 558:22]
      state <= 3'h0; // @[src/main/scala/nutcore/mem/Cache.scala 558:22]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
      if (_ismmioRec_T) begin // @[src/main/scala/nutcore/mem/Cache.scala 575:45]
        if (ismmio) begin // @[src/main/scala/nutcore/mem/Cache.scala 575:59]
          state <= 3'h3;
        end else begin
          state <= 3'h1;
        end
      end
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
      if (_T_11) begin // @[src/main/scala/nutcore/mem/Cache.scala 578:34]
        state <= 3'h2; // @[src/main/scala/nutcore/mem/Cache.scala 578:42]
      end
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
      state <= _GEN_6;
    end else begin
      state <= _GEN_12;
    end
    if (_ismmioRec_T) begin // @[src/main/scala/nutcore/mem/Cache.scala 561:28]
      ismmioRec <= ismmio; // @[src/main/scala/nutcore/mem/Cache.scala 561:28]
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/Cache.scala 570:33]
      alreadyOutFire <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 570:33]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
      alreadyOutFire <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 574:22]
    end else begin
      alreadyOutFire <= _GEN_3;
    end
    if (_ismmioRec_T) begin // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
      reqaddr <= io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    if (_ismmioRec_T) begin // @[src/main/scala/nutcore/mem/Cache.scala 595:22]
      cmd <= io_in_req_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 595:22]
    end
    if (_ismmioRec_T) begin // @[src/main/scala/nutcore/mem/Cache.scala 596:23]
      size <= io_in_req_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 596:23]
    end
    if (_ismmioRec_T) begin // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
      wdata <= io_in_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    if (_ismmioRec_T) begin // @[src/main/scala/nutcore/mem/Cache.scala 598:24]
      wmask <= io_in_req_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 598:24]
    end
    if (_T_17) begin // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
      mmiordata <= io_mmio_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    if (_T_17) begin // @[src/main/scala/nutcore/mem/Cache.scala 604:26]
      mmiocmd <= io_mmio_resp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 604:26]
    end
    if (_T_13) begin // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
      memrdata <= io_out_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    if (_T_13) begin // @[src/main/scala/nutcore/mem/Cache.scala 606:25]
      memcmd <= io_out_mem_resp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 606:25]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  ismmioRec = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  alreadyOutFire = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  reqaddr = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  cmd = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  size = _RAND_5[2:0];
  _RAND_6 = {2{`RANDOM}};
  wdata = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  wmask = _RAND_7[7:0];
  _RAND_8 = {2{`RANDOM}};
  mmiordata = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  mmiocmd = _RAND_9[3:0];
  _RAND_10 = {2{`RANDOM}};
  memrdata = _RAND_10[63:0];
  _RAND_11 = {1{`RANDOM}};
  memcmd = _RAND_11[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module NutCore(
  input         clock,
  input         reset,
  input         io_imem_mem_req_ready, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  output        io_imem_mem_req_valid, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  output [31:0] io_imem_mem_req_bits_addr, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  output [2:0]  io_imem_mem_req_bits_size, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  output [3:0]  io_imem_mem_req_bits_cmd, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  output [7:0]  io_imem_mem_req_bits_wmask, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  output [63:0] io_imem_mem_req_bits_wdata, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  output        io_imem_mem_resp_ready, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  input         io_imem_mem_resp_valid, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  input  [3:0]  io_imem_mem_resp_bits_cmd, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  input  [63:0] io_imem_mem_resp_bits_rdata, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  output        io_imem_coh_req_ready, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  input         io_imem_coh_req_valid, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  input  [31:0] io_imem_coh_req_bits_addr, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  input  [2:0]  io_imem_coh_req_bits_size, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  input  [3:0]  io_imem_coh_req_bits_cmd, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  input  [7:0]  io_imem_coh_req_bits_wmask, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  input  [63:0] io_imem_coh_req_bits_wdata, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  input         io_imem_coh_resp_ready, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  output        io_imem_coh_resp_valid, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  output [3:0]  io_imem_coh_resp_bits_cmd, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  output [63:0] io_imem_coh_resp_bits_rdata, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  input         io_dmem_mem_req_ready, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  output        io_dmem_mem_req_valid, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  output [31:0] io_dmem_mem_req_bits_addr, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  output [2:0]  io_dmem_mem_req_bits_size, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  output [3:0]  io_dmem_mem_req_bits_cmd, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  output [7:0]  io_dmem_mem_req_bits_wmask, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  output [63:0] io_dmem_mem_req_bits_wdata, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  output        io_dmem_mem_resp_ready, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  input         io_dmem_mem_resp_valid, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  input  [3:0]  io_dmem_mem_resp_bits_cmd, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  input  [63:0] io_dmem_mem_resp_bits_rdata, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  output        io_dmem_coh_req_ready, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  input         io_dmem_coh_req_valid, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  input  [31:0] io_dmem_coh_req_bits_addr, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  input  [2:0]  io_dmem_coh_req_bits_size, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  input  [3:0]  io_dmem_coh_req_bits_cmd, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  input  [7:0]  io_dmem_coh_req_bits_wmask, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  input  [63:0] io_dmem_coh_req_bits_wdata, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  input         io_dmem_coh_resp_ready, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  output        io_dmem_coh_resp_valid, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  output [3:0]  io_dmem_coh_resp_bits_cmd, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  output [63:0] io_dmem_coh_resp_bits_rdata, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  input         io_mmio_req_ready, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  output        io_mmio_req_valid, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  output [31:0] io_mmio_req_bits_addr, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  output [2:0]  io_mmio_req_bits_size, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  output [3:0]  io_mmio_req_bits_cmd, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  output [7:0]  io_mmio_req_bits_wmask, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  output [63:0] io_mmio_req_bits_wdata, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  output        io_mmio_resp_ready, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  input         io_mmio_resp_valid, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  input  [3:0]  io_mmio_resp_bits_cmd, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  input  [63:0] io_mmio_resp_bits_rdata, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  output        io_frontend_req_ready, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  input         io_frontend_req_valid, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  input  [31:0] io_frontend_req_bits_addr, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  input  [2:0]  io_frontend_req_bits_size, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  input  [3:0]  io_frontend_req_bits_cmd, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  input  [7:0]  io_frontend_req_bits_wmask, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  input  [63:0] io_frontend_req_bits_wdata, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  input         io_frontend_resp_ready, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  output        io_frontend_resp_valid, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  output [3:0]  io_frontend_resp_bits_cmd, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  output [63:0] io_frontend_resp_bits_rdata, // @[src/main/scala/nutcore/NutCore.scala 114:14]
  output        rvfi_valid, // @[src/main/scala/nutcore/NutCore.scala 115:16]
  output [63:0] rvfi_order, // @[src/main/scala/nutcore/NutCore.scala 115:16]
  output [63:0] rvfi_insn, // @[src/main/scala/nutcore/NutCore.scala 115:16]
  output        rvfi_trap, // @[src/main/scala/nutcore/NutCore.scala 115:16]
  output        rvfi_halt, // @[src/main/scala/nutcore/NutCore.scala 115:16]
  output        rvfi_intr, // @[src/main/scala/nutcore/NutCore.scala 115:16]
  output [1:0]  rvfi_mode, // @[src/main/scala/nutcore/NutCore.scala 115:16]
  output [1:0]  rvfi_ixl, // @[src/main/scala/nutcore/NutCore.scala 115:16]
  output [4:0]  rvfi_rs1_addr, // @[src/main/scala/nutcore/NutCore.scala 115:16]
  output [4:0]  rvfi_rs2_addr, // @[src/main/scala/nutcore/NutCore.scala 115:16]
  output [63:0] rvfi_rs1_rdata, // @[src/main/scala/nutcore/NutCore.scala 115:16]
  output [63:0] rvfi_rs2_rdata, // @[src/main/scala/nutcore/NutCore.scala 115:16]
  output [4:0]  rvfi_rd_addr, // @[src/main/scala/nutcore/NutCore.scala 115:16]
  output [63:0] rvfi_rd_wdata, // @[src/main/scala/nutcore/NutCore.scala 115:16]
  output [63:0] rvfi_pc_rdata, // @[src/main/scala/nutcore/NutCore.scala 115:16]
  output [63:0] rvfi_pc_wdata, // @[src/main/scala/nutcore/NutCore.scala 115:16]
  output [63:0] rvfi_mem_addr, // @[src/main/scala/nutcore/NutCore.scala 115:16]
  output [7:0]  rvfi_mem_rmask, // @[src/main/scala/nutcore/NutCore.scala 115:16]
  output [7:0]  rvfi_mem_wmask, // @[src/main/scala/nutcore/NutCore.scala 115:16]
  output [63:0] rvfi_mem_rdata, // @[src/main/scala/nutcore/NutCore.scala 115:16]
  output [63:0] rvfi_mem_wdata // @[src/main/scala/nutcore/NutCore.scala 115:16]
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [63:0] _RAND_80;
  reg [63:0] _RAND_81;
  reg [63:0] _RAND_82;
  reg [63:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [63:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
`endif // RANDOMIZE_REG_INIT
  wire  frontend_clock; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  frontend_reset; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  frontend_io_imem_req_ready; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  frontend_io_imem_req_valid; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire [38:0] frontend_io_imem_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire [86:0] frontend_io_imem_req_bits_user; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  frontend_io_imem_resp_ready; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  frontend_io_imem_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire [63:0] frontend_io_imem_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire [86:0] frontend_io_imem_resp_bits_user; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  frontend_io_out_0_ready; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  frontend_io_out_0_valid; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire [63:0] frontend_io_out_0_bits_cf_instr; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire [38:0] frontend_io_out_0_bits_cf_pc; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire [38:0] frontend_io_out_0_bits_cf_pnpc; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  frontend_io_out_0_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  frontend_io_out_0_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  frontend_io_out_0_bits_cf_intrVec_0; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  frontend_io_out_0_bits_cf_intrVec_1; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  frontend_io_out_0_bits_cf_intrVec_2; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  frontend_io_out_0_bits_cf_intrVec_3; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  frontend_io_out_0_bits_cf_intrVec_4; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  frontend_io_out_0_bits_cf_intrVec_5; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  frontend_io_out_0_bits_cf_intrVec_6; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  frontend_io_out_0_bits_cf_intrVec_7; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  frontend_io_out_0_bits_cf_intrVec_8; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  frontend_io_out_0_bits_cf_intrVec_9; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  frontend_io_out_0_bits_cf_intrVec_10; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  frontend_io_out_0_bits_cf_intrVec_11; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire [3:0] frontend_io_out_0_bits_cf_brIdx; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  frontend_io_out_0_bits_ctrl_src1Type; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  frontend_io_out_0_bits_ctrl_src2Type; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire [2:0] frontend_io_out_0_bits_ctrl_fuType; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire [6:0] frontend_io_out_0_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire [4:0] frontend_io_out_0_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire [4:0] frontend_io_out_0_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  frontend_io_out_0_bits_ctrl_rfWen; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire [4:0] frontend_io_out_0_bits_ctrl_rfDest; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire [63:0] frontend_io_out_0_bits_data_imm; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  frontend_io_out_1_bits_cf_intrVec_0; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  frontend_io_out_1_bits_cf_intrVec_1; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  frontend_io_out_1_bits_cf_intrVec_2; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  frontend_io_out_1_bits_cf_intrVec_3; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  frontend_io_out_1_bits_cf_intrVec_4; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  frontend_io_out_1_bits_cf_intrVec_5; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  frontend_io_out_1_bits_cf_intrVec_6; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  frontend_io_out_1_bits_cf_intrVec_7; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  frontend_io_out_1_bits_cf_intrVec_8; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  frontend_io_out_1_bits_cf_intrVec_9; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  frontend_io_out_1_bits_cf_intrVec_10; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  frontend_io_out_1_bits_cf_intrVec_11; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire [3:0] frontend_io_flushVec; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire [38:0] frontend_io_redirect_target; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  frontend_io_redirect_valid; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  frontend_flushICache; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  frontend_REG_valid; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire [38:0] frontend_REG_pc; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  frontend_REG_isMissPredict; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire [38:0] frontend_REG_actualTarget; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  frontend_REG_actualTaken; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire [6:0] frontend_REG_fuOpType; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire [1:0] frontend_REG_btbType; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  frontend_REG_isRVC; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire [11:0] frontend_intrVec; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  frontend_flushTLB; // @[src/main/scala/nutcore/NutCore.scala 142:34]
  wire  backend_clock; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire  backend_reset; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire  backend_io_in_0_ready; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire  backend_io_in_0_valid; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire [63:0] backend_io_in_0_bits_cf_instr; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire [38:0] backend_io_in_0_bits_cf_pc; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire [38:0] backend_io_in_0_bits_cf_pnpc; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire  backend_io_in_0_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire  backend_io_in_0_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire  backend_io_in_0_bits_cf_intrVec_0; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire  backend_io_in_0_bits_cf_intrVec_1; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire  backend_io_in_0_bits_cf_intrVec_2; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire  backend_io_in_0_bits_cf_intrVec_3; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire  backend_io_in_0_bits_cf_intrVec_4; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire  backend_io_in_0_bits_cf_intrVec_5; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire  backend_io_in_0_bits_cf_intrVec_6; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire  backend_io_in_0_bits_cf_intrVec_7; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire  backend_io_in_0_bits_cf_intrVec_8; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire  backend_io_in_0_bits_cf_intrVec_9; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire  backend_io_in_0_bits_cf_intrVec_10; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire  backend_io_in_0_bits_cf_intrVec_11; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire [3:0] backend_io_in_0_bits_cf_brIdx; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire  backend_io_in_0_bits_ctrl_src1Type; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire  backend_io_in_0_bits_ctrl_src2Type; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire [2:0] backend_io_in_0_bits_ctrl_fuType; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire [6:0] backend_io_in_0_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire [4:0] backend_io_in_0_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire [4:0] backend_io_in_0_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire  backend_io_in_0_bits_ctrl_rfWen; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire [4:0] backend_io_in_0_bits_ctrl_rfDest; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire [63:0] backend_io_in_0_bits_data_imm; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire [1:0] backend_io_flush; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire  backend_io_dmem_req_ready; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire  backend_io_dmem_req_valid; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire [38:0] backend_io_dmem_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire [2:0] backend_io_dmem_req_bits_size; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire [3:0] backend_io_dmem_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire [7:0] backend_io_dmem_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire [63:0] backend_io_dmem_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire  backend_io_dmem_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire [63:0] backend_io_dmem_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire [38:0] backend_io_redirect_target; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire  backend_io_redirect_valid; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire [63:0] backend_io_in_bits_decode_data_src1; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire  backend__T_2_0; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire  backend_io_in_valid; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire [4:0] backend_io_in_bits_decode_ctrl_rfSrc1; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire [4:0] backend_io_wb_rfDest; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire  backend_flushICache; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire [63:0] backend_rvfi_order; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire [63:0] backend_io_in_bits_mem_rvfi_addr_real; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire [4:0] backend_io_in_bits_decode_ctrl_rfSrc2; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire  backend_REG_valid; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire [38:0] backend_REG_pc; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire  backend_REG_isMissPredict; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire [38:0] backend_REG_actualTarget; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire  backend_REG_actualTaken; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire [6:0] backend_REG_fuOpType; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire [1:0] backend_REG_btbType; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire  backend_REG_isRVC; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire [63:0] backend__T_145; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire [63:0] backend_io_in_bits_mem_rvfi_rdata; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire [63:0] backend__T_151; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire [63:0] backend_io_in_bits_decode_cf_instr; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire  backend_REG_0; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire [63:0] backend_io_in_bits_mem_rvfi_wdata; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire [63:0] backend__T_142; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire [63:0] backend_io_in_bits_decode_data_src2; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire [11:0] backend_intrVec; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire [7:0] backend_io_in_bits_mem_rvfi_rmask; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire  backend_flushTLB; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire [7:0] backend_io_in_bits_mem_rvfi_wmask; // @[src/main/scala/nutcore/NutCore.scala 185:25]
  wire  mmioXbar_clock; // @[src/main/scala/nutcore/NutCore.scala 189:26]
  wire  mmioXbar_reset; // @[src/main/scala/nutcore/NutCore.scala 189:26]
  wire  mmioXbar_io_in_0_req_ready; // @[src/main/scala/nutcore/NutCore.scala 189:26]
  wire  mmioXbar_io_in_0_req_valid; // @[src/main/scala/nutcore/NutCore.scala 189:26]
  wire [31:0] mmioXbar_io_in_0_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 189:26]
  wire  mmioXbar_io_in_0_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 189:26]
  wire [63:0] mmioXbar_io_in_0_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 189:26]
  wire  mmioXbar_io_in_1_req_ready; // @[src/main/scala/nutcore/NutCore.scala 189:26]
  wire  mmioXbar_io_in_1_req_valid; // @[src/main/scala/nutcore/NutCore.scala 189:26]
  wire [31:0] mmioXbar_io_in_1_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 189:26]
  wire [2:0] mmioXbar_io_in_1_req_bits_size; // @[src/main/scala/nutcore/NutCore.scala 189:26]
  wire [3:0] mmioXbar_io_in_1_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 189:26]
  wire [7:0] mmioXbar_io_in_1_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 189:26]
  wire [63:0] mmioXbar_io_in_1_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 189:26]
  wire  mmioXbar_io_in_1_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 189:26]
  wire [3:0] mmioXbar_io_in_1_resp_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 189:26]
  wire [63:0] mmioXbar_io_in_1_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 189:26]
  wire  mmioXbar_io_out_req_ready; // @[src/main/scala/nutcore/NutCore.scala 189:26]
  wire  mmioXbar_io_out_req_valid; // @[src/main/scala/nutcore/NutCore.scala 189:26]
  wire [31:0] mmioXbar_io_out_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 189:26]
  wire [2:0] mmioXbar_io_out_req_bits_size; // @[src/main/scala/nutcore/NutCore.scala 189:26]
  wire [3:0] mmioXbar_io_out_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 189:26]
  wire [7:0] mmioXbar_io_out_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 189:26]
  wire [63:0] mmioXbar_io_out_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 189:26]
  wire  mmioXbar_io_out_resp_ready; // @[src/main/scala/nutcore/NutCore.scala 189:26]
  wire  mmioXbar_io_out_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 189:26]
  wire [3:0] mmioXbar_io_out_resp_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 189:26]
  wire [63:0] mmioXbar_io_out_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 189:26]
  wire  dmemXbar_clock; // @[src/main/scala/nutcore/NutCore.scala 190:26]
  wire  dmemXbar_reset; // @[src/main/scala/nutcore/NutCore.scala 190:26]
  wire  dmemXbar_io_in_0_req_ready; // @[src/main/scala/nutcore/NutCore.scala 190:26]
  wire  dmemXbar_io_in_0_req_valid; // @[src/main/scala/nutcore/NutCore.scala 190:26]
  wire [31:0] dmemXbar_io_in_0_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 190:26]
  wire [2:0] dmemXbar_io_in_0_req_bits_size; // @[src/main/scala/nutcore/NutCore.scala 190:26]
  wire [3:0] dmemXbar_io_in_0_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 190:26]
  wire [7:0] dmemXbar_io_in_0_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 190:26]
  wire [63:0] dmemXbar_io_in_0_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 190:26]
  wire  dmemXbar_io_in_0_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 190:26]
  wire [63:0] dmemXbar_io_in_0_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 190:26]
  wire  dmemXbar_io_in_3_req_ready; // @[src/main/scala/nutcore/NutCore.scala 190:26]
  wire  dmemXbar_io_in_3_req_valid; // @[src/main/scala/nutcore/NutCore.scala 190:26]
  wire [31:0] dmemXbar_io_in_3_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 190:26]
  wire [2:0] dmemXbar_io_in_3_req_bits_size; // @[src/main/scala/nutcore/NutCore.scala 190:26]
  wire [3:0] dmemXbar_io_in_3_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 190:26]
  wire [7:0] dmemXbar_io_in_3_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 190:26]
  wire [63:0] dmemXbar_io_in_3_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 190:26]
  wire  dmemXbar_io_in_3_resp_ready; // @[src/main/scala/nutcore/NutCore.scala 190:26]
  wire  dmemXbar_io_in_3_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 190:26]
  wire [3:0] dmemXbar_io_in_3_resp_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 190:26]
  wire [63:0] dmemXbar_io_in_3_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 190:26]
  wire  dmemXbar_io_out_req_ready; // @[src/main/scala/nutcore/NutCore.scala 190:26]
  wire  dmemXbar_io_out_req_valid; // @[src/main/scala/nutcore/NutCore.scala 190:26]
  wire [31:0] dmemXbar_io_out_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 190:26]
  wire [2:0] dmemXbar_io_out_req_bits_size; // @[src/main/scala/nutcore/NutCore.scala 190:26]
  wire [3:0] dmemXbar_io_out_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 190:26]
  wire [7:0] dmemXbar_io_out_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 190:26]
  wire [63:0] dmemXbar_io_out_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 190:26]
  wire  dmemXbar_io_out_resp_ready; // @[src/main/scala/nutcore/NutCore.scala 190:26]
  wire  dmemXbar_io_out_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 190:26]
  wire [3:0] dmemXbar_io_out_resp_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 190:26]
  wire [63:0] dmemXbar_io_out_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 190:26]
  wire  itlb_io_in_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 438:13]
  wire  itlb_io_in_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 438:13]
  wire [38:0] itlb_io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 438:13]
  wire [86:0] itlb_io_in_req_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 438:13]
  wire  itlb_io_in_resp_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 438:13]
  wire  itlb_io_in_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 438:13]
  wire [63:0] itlb_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 438:13]
  wire [86:0] itlb_io_in_resp_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 438:13]
  wire  itlb_io_out_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 438:13]
  wire  itlb_io_out_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 438:13]
  wire [31:0] itlb_io_out_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 438:13]
  wire [86:0] itlb_io_out_req_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 438:13]
  wire  itlb_io_out_resp_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 438:13]
  wire  itlb_io_out_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 438:13]
  wire [63:0] itlb_io_out_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 438:13]
  wire [86:0] itlb_io_out_resp_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 438:13]
  wire  io_imem_cache_clock; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_reset; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_in_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_in_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [31:0] io_imem_cache_io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [86:0] io_imem_cache_io_in_req_bits_user; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_in_resp_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_in_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [63:0] io_imem_cache_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [86:0] io_imem_cache_io_in_resp_bits_user; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [1:0] io_imem_cache_io_flush; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_out_mem_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_out_mem_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [31:0] io_imem_cache_io_out_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_out_mem_resp_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_out_mem_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [63:0] io_imem_cache_io_out_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_mmio_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_mmio_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [31:0] io_imem_cache_io_mmio_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_mmio_resp_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_mmio_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [63:0] io_imem_cache_io_mmio_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  dtlb_io_in_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 438:13]
  wire  dtlb_io_in_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 438:13]
  wire [38:0] dtlb_io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 438:13]
  wire [2:0] dtlb_io_in_req_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 438:13]
  wire [3:0] dtlb_io_in_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 438:13]
  wire [7:0] dtlb_io_in_req_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 438:13]
  wire [63:0] dtlb_io_in_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 438:13]
  wire  dtlb_io_in_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 438:13]
  wire [63:0] dtlb_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 438:13]
  wire  dtlb_io_out_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 438:13]
  wire  dtlb_io_out_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 438:13]
  wire [31:0] dtlb_io_out_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 438:13]
  wire [2:0] dtlb_io_out_req_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 438:13]
  wire [3:0] dtlb_io_out_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 438:13]
  wire [7:0] dtlb_io_out_req_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 438:13]
  wire [63:0] dtlb_io_out_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 438:13]
  wire  dtlb_io_out_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 438:13]
  wire [63:0] dtlb_io_out_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 438:13]
  wire  io_dmem_cache_clock; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_reset; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_in_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_in_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [31:0] io_dmem_cache_io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [2:0] io_dmem_cache_io_in_req_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [3:0] io_dmem_cache_io_in_req_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [7:0] io_dmem_cache_io_in_req_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [63:0] io_dmem_cache_io_in_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_in_resp_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_in_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [3:0] io_dmem_cache_io_in_resp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [63:0] io_dmem_cache_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_out_mem_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_out_mem_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [31:0] io_dmem_cache_io_out_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [2:0] io_dmem_cache_io_out_mem_req_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [3:0] io_dmem_cache_io_out_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [7:0] io_dmem_cache_io_out_mem_req_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [63:0] io_dmem_cache_io_out_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_out_mem_resp_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_out_mem_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [3:0] io_dmem_cache_io_out_mem_resp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [63:0] io_dmem_cache_io_out_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_mmio_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_mmio_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [31:0] io_dmem_cache_io_mmio_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [2:0] io_dmem_cache_io_mmio_req_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [3:0] io_dmem_cache_io_mmio_req_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [7:0] io_dmem_cache_io_mmio_req_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [63:0] io_dmem_cache_io_mmio_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_mmio_resp_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_mmio_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [3:0] io_dmem_cache_io_mmio_resp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [63:0] io_dmem_cache_io_mmio_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  _T_1 = ~reset; // @[src/main/scala/nutcore/NutCore.scala 132:9]
  wire  someassumeid = backend__T_2_0;
  reg [63:0] dataBuffer_0_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [38:0] dataBuffer_0_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [38:0] dataBuffer_0_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_intrVec_0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_intrVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_intrVec_4; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_intrVec_6; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_intrVec_8; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_intrVec_10; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [3:0] dataBuffer_0_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [2:0] dataBuffer_0_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [6:0] dataBuffer_0_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_0_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_0_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_0_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [63:0] dataBuffer_0_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [63:0] dataBuffer_1_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [38:0] dataBuffer_1_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [38:0] dataBuffer_1_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_intrVec_0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_intrVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_intrVec_4; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_intrVec_6; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_intrVec_8; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_intrVec_10; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [3:0] dataBuffer_1_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [2:0] dataBuffer_1_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [6:0] dataBuffer_1_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_1_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_1_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_1_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [63:0] dataBuffer_1_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [63:0] dataBuffer_2_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [38:0] dataBuffer_2_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [38:0] dataBuffer_2_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_intrVec_0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_intrVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_intrVec_4; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_intrVec_6; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_intrVec_8; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_intrVec_10; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [3:0] dataBuffer_2_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [2:0] dataBuffer_2_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [6:0] dataBuffer_2_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_2_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_2_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_2_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [63:0] dataBuffer_2_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [63:0] dataBuffer_3_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [38:0] dataBuffer_3_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [38:0] dataBuffer_3_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_intrVec_0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_intrVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_intrVec_4; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_intrVec_6; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_intrVec_8; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_intrVec_10; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [3:0] dataBuffer_3_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [2:0] dataBuffer_3_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [6:0] dataBuffer_3_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_3_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_3_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_3_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [63:0] dataBuffer_3_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [1:0] ringBufferHead; // @[src/main/scala/utils/PipelineVector.scala 30:33]
  reg [1:0] ringBufferTail; // @[src/main/scala/utils/PipelineVector.scala 31:33]
  wire [1:0] _ringBufferAllowin_T_1 = ringBufferHead + 2'h1; // @[src/main/scala/utils/PipelineVector.scala 33:63]
  wire [1:0] _ringBufferAllowin_T_4 = ringBufferHead + 2'h2; // @[src/main/scala/utils/PipelineVector.scala 33:63]
  wire  ringBufferAllowin = _ringBufferAllowin_T_1 != ringBufferTail & _ringBufferAllowin_T_4 != ringBufferTail; // @[src/main/scala/utils/PipelineVector.scala 33:124]
  wire  needEnqueue_0 = frontend_io_out_0_valid; // @[src/main/scala/utils/PipelineVector.scala 36:27 37:20]
  wire [1:0] enqueueSize = {{1'd0}, needEnqueue_0}; // @[src/main/scala/utils/PipelineVector.scala 40:44]
  wire  enqueueFire_0 = enqueueSize >= 2'h1; // @[src/main/scala/utils/PipelineVector.scala 41:53]
  wire  enqueueFire_1 = enqueueSize >= 2'h2; // @[src/main/scala/utils/PipelineVector.scala 41:53]
  wire  wen = frontend_io_out_0_ready & frontend_io_out_0_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [2:0] _T_4 = {{1'd0}, ringBufferHead}; // @[src/main/scala/utils/PipelineVector.scala 45:45]
  wire [63:0] _dataBuffer_T_cf_instr = needEnqueue_0 ? frontend_io_out_0_bits_cf_instr : 64'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [38:0] _dataBuffer_T_cf_pc = needEnqueue_0 ? frontend_io_out_0_bits_cf_pc : 39'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [38:0] _dataBuffer_T_cf_pnpc = needEnqueue_0 ? frontend_io_out_0_bits_cf_pnpc : 39'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire  _dataBuffer_T_cf_intrVec_0 = needEnqueue_0 ? frontend_io_out_0_bits_cf_intrVec_0 :
    frontend_io_out_1_bits_cf_intrVec_0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire  _dataBuffer_T_cf_intrVec_1 = needEnqueue_0 ? frontend_io_out_0_bits_cf_intrVec_1 :
    frontend_io_out_1_bits_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire  _dataBuffer_T_cf_intrVec_2 = needEnqueue_0 ? frontend_io_out_0_bits_cf_intrVec_2 :
    frontend_io_out_1_bits_cf_intrVec_2; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire  _dataBuffer_T_cf_intrVec_3 = needEnqueue_0 ? frontend_io_out_0_bits_cf_intrVec_3 :
    frontend_io_out_1_bits_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire  _dataBuffer_T_cf_intrVec_4 = needEnqueue_0 ? frontend_io_out_0_bits_cf_intrVec_4 :
    frontend_io_out_1_bits_cf_intrVec_4; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire  _dataBuffer_T_cf_intrVec_5 = needEnqueue_0 ? frontend_io_out_0_bits_cf_intrVec_5 :
    frontend_io_out_1_bits_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire  _dataBuffer_T_cf_intrVec_6 = needEnqueue_0 ? frontend_io_out_0_bits_cf_intrVec_6 :
    frontend_io_out_1_bits_cf_intrVec_6; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire  _dataBuffer_T_cf_intrVec_7 = needEnqueue_0 ? frontend_io_out_0_bits_cf_intrVec_7 :
    frontend_io_out_1_bits_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire  _dataBuffer_T_cf_intrVec_8 = needEnqueue_0 ? frontend_io_out_0_bits_cf_intrVec_8 :
    frontend_io_out_1_bits_cf_intrVec_8; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire  _dataBuffer_T_cf_intrVec_9 = needEnqueue_0 ? frontend_io_out_0_bits_cf_intrVec_9 :
    frontend_io_out_1_bits_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire  _dataBuffer_T_cf_intrVec_10 = needEnqueue_0 ? frontend_io_out_0_bits_cf_intrVec_10 :
    frontend_io_out_1_bits_cf_intrVec_10; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire  _dataBuffer_T_cf_intrVec_11 = needEnqueue_0 ? frontend_io_out_0_bits_cf_intrVec_11 :
    frontend_io_out_1_bits_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [3:0] _dataBuffer_T_cf_brIdx = needEnqueue_0 ? frontend_io_out_0_bits_cf_brIdx : 4'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire  _dataBuffer_T_ctrl_src1Type = needEnqueue_0 ? frontend_io_out_0_bits_ctrl_src1Type : 1'h1; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire  _dataBuffer_T_ctrl_src2Type = needEnqueue_0 ? frontend_io_out_0_bits_ctrl_src2Type : 1'h1; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [2:0] _dataBuffer_T_ctrl_fuType = needEnqueue_0 ? frontend_io_out_0_bits_ctrl_fuType : 3'h3; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [6:0] _dataBuffer_T_ctrl_fuOpType = needEnqueue_0 ? frontend_io_out_0_bits_ctrl_fuOpType : 7'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [4:0] _dataBuffer_T_ctrl_rfSrc1 = needEnqueue_0 ? frontend_io_out_0_bits_ctrl_rfSrc1 : 5'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [4:0] _dataBuffer_T_ctrl_rfSrc2 = needEnqueue_0 ? frontend_io_out_0_bits_ctrl_rfSrc2 : 5'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [4:0] _dataBuffer_T_ctrl_rfDest = needEnqueue_0 ? frontend_io_out_0_bits_ctrl_rfDest : 5'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [63:0] _dataBuffer_T_data_imm = needEnqueue_0 ? frontend_io_out_0_bits_data_imm : 64'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [63:0] _GEN_0 = 2'h0 == _T_4[1:0] ? _dataBuffer_T_cf_instr : dataBuffer_0_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_1 = 2'h1 == _T_4[1:0] ? _dataBuffer_T_cf_instr : dataBuffer_1_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_2 = 2'h2 == _T_4[1:0] ? _dataBuffer_T_cf_instr : dataBuffer_2_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_3 = 2'h3 == _T_4[1:0] ? _dataBuffer_T_cf_instr : dataBuffer_3_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_4 = 2'h0 == _T_4[1:0] ? _dataBuffer_T_cf_pc : dataBuffer_0_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_5 = 2'h1 == _T_4[1:0] ? _dataBuffer_T_cf_pc : dataBuffer_1_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_6 = 2'h2 == _T_4[1:0] ? _dataBuffer_T_cf_pc : dataBuffer_2_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_7 = 2'h3 == _T_4[1:0] ? _dataBuffer_T_cf_pc : dataBuffer_3_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_8 = 2'h0 == _T_4[1:0] ? _dataBuffer_T_cf_pnpc : dataBuffer_0_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_9 = 2'h1 == _T_4[1:0] ? _dataBuffer_T_cf_pnpc : dataBuffer_1_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_10 = 2'h2 == _T_4[1:0] ? _dataBuffer_T_cf_pnpc : dataBuffer_2_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_11 = 2'h3 == _T_4[1:0] ? _dataBuffer_T_cf_pnpc : dataBuffer_3_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_28 = 2'h0 == _T_4[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_1 :
    dataBuffer_0_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_29 = 2'h1 == _T_4[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_1 :
    dataBuffer_1_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_30 = 2'h2 == _T_4[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_1 :
    dataBuffer_2_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_31 = 2'h3 == _T_4[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_1 :
    dataBuffer_3_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_32 = 2'h0 == _T_4[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_2 :
    dataBuffer_0_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_33 = 2'h1 == _T_4[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_2 :
    dataBuffer_1_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_34 = 2'h2 == _T_4[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_2 :
    dataBuffer_2_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_35 = 2'h3 == _T_4[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_2 :
    dataBuffer_3_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_88 = 2'h0 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_0 : dataBuffer_0_cf_intrVec_0; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_89 = 2'h1 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_0 : dataBuffer_1_cf_intrVec_0; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_90 = 2'h2 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_0 : dataBuffer_2_cf_intrVec_0; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_91 = 2'h3 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_0 : dataBuffer_3_cf_intrVec_0; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_92 = 2'h0 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_1 : dataBuffer_0_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_93 = 2'h1 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_1 : dataBuffer_1_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_94 = 2'h2 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_1 : dataBuffer_2_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_95 = 2'h3 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_1 : dataBuffer_3_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_96 = 2'h0 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_2 : dataBuffer_0_cf_intrVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_97 = 2'h1 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_2 : dataBuffer_1_cf_intrVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_98 = 2'h2 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_2 : dataBuffer_2_cf_intrVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_99 = 2'h3 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_2 : dataBuffer_3_cf_intrVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_100 = 2'h0 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_3 : dataBuffer_0_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_101 = 2'h1 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_3 : dataBuffer_1_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_102 = 2'h2 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_3 : dataBuffer_2_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_103 = 2'h3 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_3 : dataBuffer_3_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_104 = 2'h0 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_4 : dataBuffer_0_cf_intrVec_4; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_105 = 2'h1 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_4 : dataBuffer_1_cf_intrVec_4; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_106 = 2'h2 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_4 : dataBuffer_2_cf_intrVec_4; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_107 = 2'h3 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_4 : dataBuffer_3_cf_intrVec_4; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_108 = 2'h0 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_5 : dataBuffer_0_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_109 = 2'h1 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_5 : dataBuffer_1_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_110 = 2'h2 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_5 : dataBuffer_2_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_111 = 2'h3 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_5 : dataBuffer_3_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_112 = 2'h0 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_6 : dataBuffer_0_cf_intrVec_6; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_113 = 2'h1 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_6 : dataBuffer_1_cf_intrVec_6; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_114 = 2'h2 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_6 : dataBuffer_2_cf_intrVec_6; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_115 = 2'h3 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_6 : dataBuffer_3_cf_intrVec_6; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_116 = 2'h0 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_7 : dataBuffer_0_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_117 = 2'h1 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_7 : dataBuffer_1_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_118 = 2'h2 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_7 : dataBuffer_2_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_119 = 2'h3 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_7 : dataBuffer_3_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_120 = 2'h0 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_8 : dataBuffer_0_cf_intrVec_8; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_121 = 2'h1 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_8 : dataBuffer_1_cf_intrVec_8; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_122 = 2'h2 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_8 : dataBuffer_2_cf_intrVec_8; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_123 = 2'h3 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_8 : dataBuffer_3_cf_intrVec_8; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_124 = 2'h0 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_9 : dataBuffer_0_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_125 = 2'h1 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_9 : dataBuffer_1_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_126 = 2'h2 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_9 : dataBuffer_2_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_127 = 2'h3 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_9 : dataBuffer_3_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_128 = 2'h0 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_10 : dataBuffer_0_cf_intrVec_10; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_129 = 2'h1 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_10 : dataBuffer_1_cf_intrVec_10; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_130 = 2'h2 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_10 : dataBuffer_2_cf_intrVec_10; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_131 = 2'h3 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_10 : dataBuffer_3_cf_intrVec_10; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_132 = 2'h0 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_11 : dataBuffer_0_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_133 = 2'h1 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_11 : dataBuffer_1_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_134 = 2'h2 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_11 : dataBuffer_2_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_135 = 2'h3 == _T_4[1:0] ? _dataBuffer_T_cf_intrVec_11 : dataBuffer_3_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [3:0] _GEN_136 = 2'h0 == _T_4[1:0] ? _dataBuffer_T_cf_brIdx : dataBuffer_0_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [3:0] _GEN_137 = 2'h1 == _T_4[1:0] ? _dataBuffer_T_cf_brIdx : dataBuffer_1_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [3:0] _GEN_138 = 2'h2 == _T_4[1:0] ? _dataBuffer_T_cf_brIdx : dataBuffer_2_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [3:0] _GEN_139 = 2'h3 == _T_4[1:0] ? _dataBuffer_T_cf_brIdx : dataBuffer_3_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_156 = 2'h0 == _T_4[1:0] ? _dataBuffer_T_ctrl_src1Type : dataBuffer_0_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_157 = 2'h1 == _T_4[1:0] ? _dataBuffer_T_ctrl_src1Type : dataBuffer_1_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_158 = 2'h2 == _T_4[1:0] ? _dataBuffer_T_ctrl_src1Type : dataBuffer_2_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_159 = 2'h3 == _T_4[1:0] ? _dataBuffer_T_ctrl_src1Type : dataBuffer_3_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_160 = 2'h0 == _T_4[1:0] ? _dataBuffer_T_ctrl_src2Type : dataBuffer_0_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_161 = 2'h1 == _T_4[1:0] ? _dataBuffer_T_ctrl_src2Type : dataBuffer_1_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_162 = 2'h2 == _T_4[1:0] ? _dataBuffer_T_ctrl_src2Type : dataBuffer_2_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_163 = 2'h3 == _T_4[1:0] ? _dataBuffer_T_ctrl_src2Type : dataBuffer_3_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [2:0] _GEN_164 = 2'h0 == _T_4[1:0] ? _dataBuffer_T_ctrl_fuType : dataBuffer_0_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [2:0] _GEN_165 = 2'h1 == _T_4[1:0] ? _dataBuffer_T_ctrl_fuType : dataBuffer_1_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [2:0] _GEN_166 = 2'h2 == _T_4[1:0] ? _dataBuffer_T_ctrl_fuType : dataBuffer_2_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [2:0] _GEN_167 = 2'h3 == _T_4[1:0] ? _dataBuffer_T_ctrl_fuType : dataBuffer_3_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [6:0] _GEN_168 = 2'h0 == _T_4[1:0] ? _dataBuffer_T_ctrl_fuOpType : dataBuffer_0_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [6:0] _GEN_169 = 2'h1 == _T_4[1:0] ? _dataBuffer_T_ctrl_fuOpType : dataBuffer_1_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [6:0] _GEN_170 = 2'h2 == _T_4[1:0] ? _dataBuffer_T_ctrl_fuOpType : dataBuffer_2_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [6:0] _GEN_171 = 2'h3 == _T_4[1:0] ? _dataBuffer_T_ctrl_fuOpType : dataBuffer_3_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_172 = 2'h0 == _T_4[1:0] ? _dataBuffer_T_ctrl_rfSrc1 : dataBuffer_0_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_173 = 2'h1 == _T_4[1:0] ? _dataBuffer_T_ctrl_rfSrc1 : dataBuffer_1_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_174 = 2'h2 == _T_4[1:0] ? _dataBuffer_T_ctrl_rfSrc1 : dataBuffer_2_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_175 = 2'h3 == _T_4[1:0] ? _dataBuffer_T_ctrl_rfSrc1 : dataBuffer_3_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_176 = 2'h0 == _T_4[1:0] ? _dataBuffer_T_ctrl_rfSrc2 : dataBuffer_0_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_177 = 2'h1 == _T_4[1:0] ? _dataBuffer_T_ctrl_rfSrc2 : dataBuffer_1_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_178 = 2'h2 == _T_4[1:0] ? _dataBuffer_T_ctrl_rfSrc2 : dataBuffer_2_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_179 = 2'h3 == _T_4[1:0] ? _dataBuffer_T_ctrl_rfSrc2 : dataBuffer_3_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_180 = 2'h0 == _T_4[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_rfWen : dataBuffer_0_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_181 = 2'h1 == _T_4[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_rfWen : dataBuffer_1_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_182 = 2'h2 == _T_4[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_rfWen : dataBuffer_2_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_183 = 2'h3 == _T_4[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_rfWen : dataBuffer_3_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_184 = 2'h0 == _T_4[1:0] ? _dataBuffer_T_ctrl_rfDest : dataBuffer_0_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_185 = 2'h1 == _T_4[1:0] ? _dataBuffer_T_ctrl_rfDest : dataBuffer_1_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_186 = 2'h2 == _T_4[1:0] ? _dataBuffer_T_ctrl_rfDest : dataBuffer_2_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_187 = 2'h3 == _T_4[1:0] ? _dataBuffer_T_ctrl_rfDest : dataBuffer_3_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_216 = 2'h0 == _T_4[1:0] ? _dataBuffer_T_data_imm : dataBuffer_0_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_217 = 2'h1 == _T_4[1:0] ? _dataBuffer_T_data_imm : dataBuffer_1_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_218 = 2'h2 == _T_4[1:0] ? _dataBuffer_T_data_imm : dataBuffer_2_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_219 = 2'h3 == _T_4[1:0] ? _dataBuffer_T_data_imm : dataBuffer_3_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_220 = enqueueFire_0 ? _GEN_0 : dataBuffer_0_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_221 = enqueueFire_0 ? _GEN_1 : dataBuffer_1_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_222 = enqueueFire_0 ? _GEN_2 : dataBuffer_2_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_223 = enqueueFire_0 ? _GEN_3 : dataBuffer_3_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_224 = enqueueFire_0 ? _GEN_4 : dataBuffer_0_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_225 = enqueueFire_0 ? _GEN_5 : dataBuffer_1_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_226 = enqueueFire_0 ? _GEN_6 : dataBuffer_2_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_227 = enqueueFire_0 ? _GEN_7 : dataBuffer_3_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_228 = enqueueFire_0 ? _GEN_8 : dataBuffer_0_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_229 = enqueueFire_0 ? _GEN_9 : dataBuffer_1_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_230 = enqueueFire_0 ? _GEN_10 : dataBuffer_2_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_231 = enqueueFire_0 ? _GEN_11 : dataBuffer_3_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_248 = enqueueFire_0 ? _GEN_28 : dataBuffer_0_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_249 = enqueueFire_0 ? _GEN_29 : dataBuffer_1_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_250 = enqueueFire_0 ? _GEN_30 : dataBuffer_2_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_251 = enqueueFire_0 ? _GEN_31 : dataBuffer_3_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_252 = enqueueFire_0 ? _GEN_32 : dataBuffer_0_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_253 = enqueueFire_0 ? _GEN_33 : dataBuffer_1_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_254 = enqueueFire_0 ? _GEN_34 : dataBuffer_2_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_255 = enqueueFire_0 ? _GEN_35 : dataBuffer_3_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_308 = enqueueFire_0 ? _GEN_88 : dataBuffer_0_cf_intrVec_0; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_309 = enqueueFire_0 ? _GEN_89 : dataBuffer_1_cf_intrVec_0; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_310 = enqueueFire_0 ? _GEN_90 : dataBuffer_2_cf_intrVec_0; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_311 = enqueueFire_0 ? _GEN_91 : dataBuffer_3_cf_intrVec_0; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_312 = enqueueFire_0 ? _GEN_92 : dataBuffer_0_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_313 = enqueueFire_0 ? _GEN_93 : dataBuffer_1_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_314 = enqueueFire_0 ? _GEN_94 : dataBuffer_2_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_315 = enqueueFire_0 ? _GEN_95 : dataBuffer_3_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_316 = enqueueFire_0 ? _GEN_96 : dataBuffer_0_cf_intrVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_317 = enqueueFire_0 ? _GEN_97 : dataBuffer_1_cf_intrVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_318 = enqueueFire_0 ? _GEN_98 : dataBuffer_2_cf_intrVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_319 = enqueueFire_0 ? _GEN_99 : dataBuffer_3_cf_intrVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_320 = enqueueFire_0 ? _GEN_100 : dataBuffer_0_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_321 = enqueueFire_0 ? _GEN_101 : dataBuffer_1_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_322 = enqueueFire_0 ? _GEN_102 : dataBuffer_2_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_323 = enqueueFire_0 ? _GEN_103 : dataBuffer_3_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_324 = enqueueFire_0 ? _GEN_104 : dataBuffer_0_cf_intrVec_4; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_325 = enqueueFire_0 ? _GEN_105 : dataBuffer_1_cf_intrVec_4; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_326 = enqueueFire_0 ? _GEN_106 : dataBuffer_2_cf_intrVec_4; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_327 = enqueueFire_0 ? _GEN_107 : dataBuffer_3_cf_intrVec_4; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_328 = enqueueFire_0 ? _GEN_108 : dataBuffer_0_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_329 = enqueueFire_0 ? _GEN_109 : dataBuffer_1_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_330 = enqueueFire_0 ? _GEN_110 : dataBuffer_2_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_331 = enqueueFire_0 ? _GEN_111 : dataBuffer_3_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_332 = enqueueFire_0 ? _GEN_112 : dataBuffer_0_cf_intrVec_6; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_333 = enqueueFire_0 ? _GEN_113 : dataBuffer_1_cf_intrVec_6; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_334 = enqueueFire_0 ? _GEN_114 : dataBuffer_2_cf_intrVec_6; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_335 = enqueueFire_0 ? _GEN_115 : dataBuffer_3_cf_intrVec_6; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_336 = enqueueFire_0 ? _GEN_116 : dataBuffer_0_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_337 = enqueueFire_0 ? _GEN_117 : dataBuffer_1_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_338 = enqueueFire_0 ? _GEN_118 : dataBuffer_2_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_339 = enqueueFire_0 ? _GEN_119 : dataBuffer_3_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_340 = enqueueFire_0 ? _GEN_120 : dataBuffer_0_cf_intrVec_8; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_341 = enqueueFire_0 ? _GEN_121 : dataBuffer_1_cf_intrVec_8; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_342 = enqueueFire_0 ? _GEN_122 : dataBuffer_2_cf_intrVec_8; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_343 = enqueueFire_0 ? _GEN_123 : dataBuffer_3_cf_intrVec_8; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_344 = enqueueFire_0 ? _GEN_124 : dataBuffer_0_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_345 = enqueueFire_0 ? _GEN_125 : dataBuffer_1_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_346 = enqueueFire_0 ? _GEN_126 : dataBuffer_2_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_347 = enqueueFire_0 ? _GEN_127 : dataBuffer_3_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_348 = enqueueFire_0 ? _GEN_128 : dataBuffer_0_cf_intrVec_10; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_349 = enqueueFire_0 ? _GEN_129 : dataBuffer_1_cf_intrVec_10; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_350 = enqueueFire_0 ? _GEN_130 : dataBuffer_2_cf_intrVec_10; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_351 = enqueueFire_0 ? _GEN_131 : dataBuffer_3_cf_intrVec_10; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_352 = enqueueFire_0 ? _GEN_132 : dataBuffer_0_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_353 = enqueueFire_0 ? _GEN_133 : dataBuffer_1_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_354 = enqueueFire_0 ? _GEN_134 : dataBuffer_2_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_355 = enqueueFire_0 ? _GEN_135 : dataBuffer_3_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_356 = enqueueFire_0 ? _GEN_136 : dataBuffer_0_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_357 = enqueueFire_0 ? _GEN_137 : dataBuffer_1_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_358 = enqueueFire_0 ? _GEN_138 : dataBuffer_2_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_359 = enqueueFire_0 ? _GEN_139 : dataBuffer_3_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_376 = enqueueFire_0 ? _GEN_156 : dataBuffer_0_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_377 = enqueueFire_0 ? _GEN_157 : dataBuffer_1_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_378 = enqueueFire_0 ? _GEN_158 : dataBuffer_2_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_379 = enqueueFire_0 ? _GEN_159 : dataBuffer_3_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_380 = enqueueFire_0 ? _GEN_160 : dataBuffer_0_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_381 = enqueueFire_0 ? _GEN_161 : dataBuffer_1_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_382 = enqueueFire_0 ? _GEN_162 : dataBuffer_2_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_383 = enqueueFire_0 ? _GEN_163 : dataBuffer_3_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [2:0] _GEN_384 = enqueueFire_0 ? _GEN_164 : dataBuffer_0_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [2:0] _GEN_385 = enqueueFire_0 ? _GEN_165 : dataBuffer_1_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [2:0] _GEN_386 = enqueueFire_0 ? _GEN_166 : dataBuffer_2_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [2:0] _GEN_387 = enqueueFire_0 ? _GEN_167 : dataBuffer_3_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [6:0] _GEN_388 = enqueueFire_0 ? _GEN_168 : dataBuffer_0_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [6:0] _GEN_389 = enqueueFire_0 ? _GEN_169 : dataBuffer_1_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [6:0] _GEN_390 = enqueueFire_0 ? _GEN_170 : dataBuffer_2_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [6:0] _GEN_391 = enqueueFire_0 ? _GEN_171 : dataBuffer_3_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_392 = enqueueFire_0 ? _GEN_172 : dataBuffer_0_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_393 = enqueueFire_0 ? _GEN_173 : dataBuffer_1_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_394 = enqueueFire_0 ? _GEN_174 : dataBuffer_2_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_395 = enqueueFire_0 ? _GEN_175 : dataBuffer_3_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_396 = enqueueFire_0 ? _GEN_176 : dataBuffer_0_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_397 = enqueueFire_0 ? _GEN_177 : dataBuffer_1_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_398 = enqueueFire_0 ? _GEN_178 : dataBuffer_2_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_399 = enqueueFire_0 ? _GEN_179 : dataBuffer_3_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_400 = enqueueFire_0 ? _GEN_180 : dataBuffer_0_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_401 = enqueueFire_0 ? _GEN_181 : dataBuffer_1_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_402 = enqueueFire_0 ? _GEN_182 : dataBuffer_2_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_403 = enqueueFire_0 ? _GEN_183 : dataBuffer_3_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_404 = enqueueFire_0 ? _GEN_184 : dataBuffer_0_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_405 = enqueueFire_0 ? _GEN_185 : dataBuffer_1_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_406 = enqueueFire_0 ? _GEN_186 : dataBuffer_2_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_407 = enqueueFire_0 ? _GEN_187 : dataBuffer_3_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_436 = enqueueFire_0 ? _GEN_216 : dataBuffer_0_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_437 = enqueueFire_0 ? _GEN_217 : dataBuffer_1_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_438 = enqueueFire_0 ? _GEN_218 : dataBuffer_2_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_439 = enqueueFire_0 ? _GEN_219 : dataBuffer_3_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [1:0] _T_7 = 2'h1 + ringBufferHead; // @[src/main/scala/utils/PipelineVector.scala 46:45]
  wire [1:0] _ringBufferHead_T_1 = ringBufferHead + enqueueSize; // @[src/main/scala/utils/PipelineVector.scala 47:42]
  wire [63:0] _GEN_1102 = 2'h1 == ringBufferTail ? dataBuffer_1_data_imm : dataBuffer_0_data_imm; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [63:0] _GEN_1103 = 2'h2 == ringBufferTail ? dataBuffer_2_data_imm : _GEN_1102; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_1134 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_rfDest : dataBuffer_0_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_1135 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_rfDest : _GEN_1134; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1138 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_rfWen : dataBuffer_0_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1139 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_rfWen : _GEN_1138; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_1142 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_rfSrc2 : dataBuffer_0_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_1143 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_rfSrc2 : _GEN_1142; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_1146 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_rfSrc1 : dataBuffer_0_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_1147 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_rfSrc1 : _GEN_1146; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [6:0] _GEN_1150 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_fuOpType : dataBuffer_0_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [6:0] _GEN_1151 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_fuOpType : _GEN_1150; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [2:0] _GEN_1154 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_fuType : dataBuffer_0_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [2:0] _GEN_1155 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_fuType : _GEN_1154; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1158 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_src2Type : dataBuffer_0_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1159 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_src2Type : _GEN_1158; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1162 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_src1Type : dataBuffer_0_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1163 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_src1Type : _GEN_1162; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [3:0] _GEN_1182 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_brIdx : dataBuffer_0_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [3:0] _GEN_1183 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_brIdx : _GEN_1182; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1186 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_intrVec_0 : dataBuffer_0_cf_intrVec_0; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1187 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_intrVec_0 : _GEN_1186; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1190 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_intrVec_1 : dataBuffer_0_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1191 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_intrVec_1 : _GEN_1190; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1194 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_intrVec_2 : dataBuffer_0_cf_intrVec_2; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1195 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_intrVec_2 : _GEN_1194; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1198 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_intrVec_3 : dataBuffer_0_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1199 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_intrVec_3 : _GEN_1198; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1202 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_intrVec_4 : dataBuffer_0_cf_intrVec_4; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1203 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_intrVec_4 : _GEN_1202; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1206 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_intrVec_5 : dataBuffer_0_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1207 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_intrVec_5 : _GEN_1206; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1210 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_intrVec_6 : dataBuffer_0_cf_intrVec_6; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1211 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_intrVec_6 : _GEN_1210; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1214 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_intrVec_7 : dataBuffer_0_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1215 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_intrVec_7 : _GEN_1214; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1218 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_intrVec_8 : dataBuffer_0_cf_intrVec_8; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1219 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_intrVec_8 : _GEN_1218; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1222 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_intrVec_9 : dataBuffer_0_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1223 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_intrVec_9 : _GEN_1222; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1226 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_intrVec_10 : dataBuffer_0_cf_intrVec_10; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1227 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_intrVec_10 : _GEN_1226; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1230 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_intrVec_11 : dataBuffer_0_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1231 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_intrVec_11 : _GEN_1230; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1238 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_exceptionVec_1 : dataBuffer_0_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1239 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_exceptionVec_1 : _GEN_1238; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1242 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_exceptionVec_2 : dataBuffer_0_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1243 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_exceptionVec_2 : _GEN_1242; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [38:0] _GEN_1310 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_pnpc : dataBuffer_0_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [38:0] _GEN_1311 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_pnpc : _GEN_1310; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [38:0] _GEN_1314 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_pc : dataBuffer_0_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [38:0] _GEN_1315 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_pc : _GEN_1314; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [63:0] _GEN_1318 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_instr : dataBuffer_0_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [63:0] _GEN_1319 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_instr : _GEN_1318; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _dequeueSize_T = backend_io_in_0_ready & backend_io_in_0_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 52:35]
  wire [1:0] dequeueSize = {{1'd0}, _dequeueSize_T}; // @[src/main/scala/utils/PipelineVector.scala 64:40]
  wire  dequeueFire = dequeueSize > 2'h0; // @[src/main/scala/utils/PipelineVector.scala 65:35]
  wire [1:0] _ringBufferTail_T_1 = ringBufferTail + dequeueSize; // @[src/main/scala/utils/PipelineVector.scala 67:42]
  wire [63:0] rvfi_mem_addr_real = backend_io_in_bits_mem_rvfi_addr_real;
  wire [38:0] _rvfi_mem_addr_T_2 = {rvfi_mem_addr_real[38:3], 3'h0}; // @[src/main/scala/nutcore/NutCore.scala 231:59]
  wire  rvfi_mem_addr_signBit = _rvfi_mem_addr_T_2[38]; // @[src/main/scala/utils/BitUtils.scala 39:20]
  wire [24:0] _rvfi_mem_addr_T_4 = rvfi_mem_addr_signBit ? 25'h1ffffff : 25'h0; // @[src/main/scala/utils/BitUtils.scala 40:46]
  reg [31:0] pcOld; // @[src/main/scala/nutcore/NutCore.scala 255:26]
  wire [63:0] _GEN_1544 = rvfi_valid ? rvfi_pc_rdata : {{32'd0}, pcOld}; // @[src/main/scala/nutcore/NutCore.scala 256:23 257:15 255:26]
  wire [63:0] _GEN_1555 = {{32'd0}, pcOld}; // @[src/main/scala/nutcore/NutCore.scala 260:31]
  wire  _T_19 = ~rvfi_valid | _GEN_1555 != rvfi_pc_rdata; // @[src/main/scala/nutcore/NutCore.scala 260:21]
  wire [63:0] _GEN_1556 = reset ? 64'h0 : _GEN_1544; // @[src/main/scala/nutcore/NutCore.scala 255:{26,26}]
  Frontend_inorder frontend ( // @[src/main/scala/nutcore/NutCore.scala 142:34]
    .clock(frontend_clock),
    .reset(frontend_reset),
    .io_imem_req_ready(frontend_io_imem_req_ready),
    .io_imem_req_valid(frontend_io_imem_req_valid),
    .io_imem_req_bits_addr(frontend_io_imem_req_bits_addr),
    .io_imem_req_bits_user(frontend_io_imem_req_bits_user),
    .io_imem_resp_ready(frontend_io_imem_resp_ready),
    .io_imem_resp_valid(frontend_io_imem_resp_valid),
    .io_imem_resp_bits_rdata(frontend_io_imem_resp_bits_rdata),
    .io_imem_resp_bits_user(frontend_io_imem_resp_bits_user),
    .io_out_0_ready(frontend_io_out_0_ready),
    .io_out_0_valid(frontend_io_out_0_valid),
    .io_out_0_bits_cf_instr(frontend_io_out_0_bits_cf_instr),
    .io_out_0_bits_cf_pc(frontend_io_out_0_bits_cf_pc),
    .io_out_0_bits_cf_pnpc(frontend_io_out_0_bits_cf_pnpc),
    .io_out_0_bits_cf_exceptionVec_1(frontend_io_out_0_bits_cf_exceptionVec_1),
    .io_out_0_bits_cf_exceptionVec_2(frontend_io_out_0_bits_cf_exceptionVec_2),
    .io_out_0_bits_cf_intrVec_0(frontend_io_out_0_bits_cf_intrVec_0),
    .io_out_0_bits_cf_intrVec_1(frontend_io_out_0_bits_cf_intrVec_1),
    .io_out_0_bits_cf_intrVec_2(frontend_io_out_0_bits_cf_intrVec_2),
    .io_out_0_bits_cf_intrVec_3(frontend_io_out_0_bits_cf_intrVec_3),
    .io_out_0_bits_cf_intrVec_4(frontend_io_out_0_bits_cf_intrVec_4),
    .io_out_0_bits_cf_intrVec_5(frontend_io_out_0_bits_cf_intrVec_5),
    .io_out_0_bits_cf_intrVec_6(frontend_io_out_0_bits_cf_intrVec_6),
    .io_out_0_bits_cf_intrVec_7(frontend_io_out_0_bits_cf_intrVec_7),
    .io_out_0_bits_cf_intrVec_8(frontend_io_out_0_bits_cf_intrVec_8),
    .io_out_0_bits_cf_intrVec_9(frontend_io_out_0_bits_cf_intrVec_9),
    .io_out_0_bits_cf_intrVec_10(frontend_io_out_0_bits_cf_intrVec_10),
    .io_out_0_bits_cf_intrVec_11(frontend_io_out_0_bits_cf_intrVec_11),
    .io_out_0_bits_cf_brIdx(frontend_io_out_0_bits_cf_brIdx),
    .io_out_0_bits_ctrl_src1Type(frontend_io_out_0_bits_ctrl_src1Type),
    .io_out_0_bits_ctrl_src2Type(frontend_io_out_0_bits_ctrl_src2Type),
    .io_out_0_bits_ctrl_fuType(frontend_io_out_0_bits_ctrl_fuType),
    .io_out_0_bits_ctrl_fuOpType(frontend_io_out_0_bits_ctrl_fuOpType),
    .io_out_0_bits_ctrl_rfSrc1(frontend_io_out_0_bits_ctrl_rfSrc1),
    .io_out_0_bits_ctrl_rfSrc2(frontend_io_out_0_bits_ctrl_rfSrc2),
    .io_out_0_bits_ctrl_rfWen(frontend_io_out_0_bits_ctrl_rfWen),
    .io_out_0_bits_ctrl_rfDest(frontend_io_out_0_bits_ctrl_rfDest),
    .io_out_0_bits_data_imm(frontend_io_out_0_bits_data_imm),
    .io_out_1_bits_cf_intrVec_0(frontend_io_out_1_bits_cf_intrVec_0),
    .io_out_1_bits_cf_intrVec_1(frontend_io_out_1_bits_cf_intrVec_1),
    .io_out_1_bits_cf_intrVec_2(frontend_io_out_1_bits_cf_intrVec_2),
    .io_out_1_bits_cf_intrVec_3(frontend_io_out_1_bits_cf_intrVec_3),
    .io_out_1_bits_cf_intrVec_4(frontend_io_out_1_bits_cf_intrVec_4),
    .io_out_1_bits_cf_intrVec_5(frontend_io_out_1_bits_cf_intrVec_5),
    .io_out_1_bits_cf_intrVec_6(frontend_io_out_1_bits_cf_intrVec_6),
    .io_out_1_bits_cf_intrVec_7(frontend_io_out_1_bits_cf_intrVec_7),
    .io_out_1_bits_cf_intrVec_8(frontend_io_out_1_bits_cf_intrVec_8),
    .io_out_1_bits_cf_intrVec_9(frontend_io_out_1_bits_cf_intrVec_9),
    .io_out_1_bits_cf_intrVec_10(frontend_io_out_1_bits_cf_intrVec_10),
    .io_out_1_bits_cf_intrVec_11(frontend_io_out_1_bits_cf_intrVec_11),
    .io_flushVec(frontend_io_flushVec),
    .io_redirect_target(frontend_io_redirect_target),
    .io_redirect_valid(frontend_io_redirect_valid),
    .flushICache(frontend_flushICache),
    .REG_valid(frontend_REG_valid),
    .REG_pc(frontend_REG_pc),
    .REG_isMissPredict(frontend_REG_isMissPredict),
    .REG_actualTarget(frontend_REG_actualTarget),
    .REG_actualTaken(frontend_REG_actualTaken),
    .REG_fuOpType(frontend_REG_fuOpType),
    .REG_btbType(frontend_REG_btbType),
    .REG_isRVC(frontend_REG_isRVC),
    .intrVec(frontend_intrVec),
    .flushTLB(frontend_flushTLB)
  );
  Backend_inorder backend ( // @[src/main/scala/nutcore/NutCore.scala 185:25]
    .clock(backend_clock),
    .reset(backend_reset),
    .io_in_0_ready(backend_io_in_0_ready),
    .io_in_0_valid(backend_io_in_0_valid),
    .io_in_0_bits_cf_instr(backend_io_in_0_bits_cf_instr),
    .io_in_0_bits_cf_pc(backend_io_in_0_bits_cf_pc),
    .io_in_0_bits_cf_pnpc(backend_io_in_0_bits_cf_pnpc),
    .io_in_0_bits_cf_exceptionVec_1(backend_io_in_0_bits_cf_exceptionVec_1),
    .io_in_0_bits_cf_exceptionVec_2(backend_io_in_0_bits_cf_exceptionVec_2),
    .io_in_0_bits_cf_intrVec_0(backend_io_in_0_bits_cf_intrVec_0),
    .io_in_0_bits_cf_intrVec_1(backend_io_in_0_bits_cf_intrVec_1),
    .io_in_0_bits_cf_intrVec_2(backend_io_in_0_bits_cf_intrVec_2),
    .io_in_0_bits_cf_intrVec_3(backend_io_in_0_bits_cf_intrVec_3),
    .io_in_0_bits_cf_intrVec_4(backend_io_in_0_bits_cf_intrVec_4),
    .io_in_0_bits_cf_intrVec_5(backend_io_in_0_bits_cf_intrVec_5),
    .io_in_0_bits_cf_intrVec_6(backend_io_in_0_bits_cf_intrVec_6),
    .io_in_0_bits_cf_intrVec_7(backend_io_in_0_bits_cf_intrVec_7),
    .io_in_0_bits_cf_intrVec_8(backend_io_in_0_bits_cf_intrVec_8),
    .io_in_0_bits_cf_intrVec_9(backend_io_in_0_bits_cf_intrVec_9),
    .io_in_0_bits_cf_intrVec_10(backend_io_in_0_bits_cf_intrVec_10),
    .io_in_0_bits_cf_intrVec_11(backend_io_in_0_bits_cf_intrVec_11),
    .io_in_0_bits_cf_brIdx(backend_io_in_0_bits_cf_brIdx),
    .io_in_0_bits_ctrl_src1Type(backend_io_in_0_bits_ctrl_src1Type),
    .io_in_0_bits_ctrl_src2Type(backend_io_in_0_bits_ctrl_src2Type),
    .io_in_0_bits_ctrl_fuType(backend_io_in_0_bits_ctrl_fuType),
    .io_in_0_bits_ctrl_fuOpType(backend_io_in_0_bits_ctrl_fuOpType),
    .io_in_0_bits_ctrl_rfSrc1(backend_io_in_0_bits_ctrl_rfSrc1),
    .io_in_0_bits_ctrl_rfSrc2(backend_io_in_0_bits_ctrl_rfSrc2),
    .io_in_0_bits_ctrl_rfWen(backend_io_in_0_bits_ctrl_rfWen),
    .io_in_0_bits_ctrl_rfDest(backend_io_in_0_bits_ctrl_rfDest),
    .io_in_0_bits_data_imm(backend_io_in_0_bits_data_imm),
    .io_flush(backend_io_flush),
    .io_dmem_req_ready(backend_io_dmem_req_ready),
    .io_dmem_req_valid(backend_io_dmem_req_valid),
    .io_dmem_req_bits_addr(backend_io_dmem_req_bits_addr),
    .io_dmem_req_bits_size(backend_io_dmem_req_bits_size),
    .io_dmem_req_bits_cmd(backend_io_dmem_req_bits_cmd),
    .io_dmem_req_bits_wmask(backend_io_dmem_req_bits_wmask),
    .io_dmem_req_bits_wdata(backend_io_dmem_req_bits_wdata),
    .io_dmem_resp_valid(backend_io_dmem_resp_valid),
    .io_dmem_resp_bits_rdata(backend_io_dmem_resp_bits_rdata),
    .io_redirect_target(backend_io_redirect_target),
    .io_redirect_valid(backend_io_redirect_valid),
    .io_in_bits_decode_data_src1(backend_io_in_bits_decode_data_src1),
    ._T_2_0(backend__T_2_0),
    .io_in_valid(backend_io_in_valid),
    .io_in_bits_decode_ctrl_rfSrc1(backend_io_in_bits_decode_ctrl_rfSrc1),
    .io_wb_rfDest(backend_io_wb_rfDest),
    .flushICache(backend_flushICache),
    .rvfi_order(backend_rvfi_order),
    .io_in_bits_mem_rvfi_addr_real(backend_io_in_bits_mem_rvfi_addr_real),
    .io_in_bits_decode_ctrl_rfSrc2(backend_io_in_bits_decode_ctrl_rfSrc2),
    .REG_valid(backend_REG_valid),
    .REG_pc(backend_REG_pc),
    .REG_isMissPredict(backend_REG_isMissPredict),
    .REG_actualTarget(backend_REG_actualTarget),
    .REG_actualTaken(backend_REG_actualTaken),
    .REG_fuOpType(backend_REG_fuOpType),
    .REG_btbType(backend_REG_btbType),
    .REG_isRVC(backend_REG_isRVC),
    ._T_145(backend__T_145),
    .io_in_bits_mem_rvfi_rdata(backend_io_in_bits_mem_rvfi_rdata),
    ._T_151(backend__T_151),
    .io_in_bits_decode_cf_instr(backend_io_in_bits_decode_cf_instr),
    .REG_0(backend_REG_0),
    .io_in_bits_mem_rvfi_wdata(backend_io_in_bits_mem_rvfi_wdata),
    ._T_142(backend__T_142),
    .io_in_bits_decode_data_src2(backend_io_in_bits_decode_data_src2),
    .intrVec(backend_intrVec),
    .io_in_bits_mem_rvfi_rmask(backend_io_in_bits_mem_rvfi_rmask),
    .flushTLB(backend_flushTLB),
    .io_in_bits_mem_rvfi_wmask(backend_io_in_bits_mem_rvfi_wmask)
  );
  SimpleBusCrossbarNto1 mmioXbar ( // @[src/main/scala/nutcore/NutCore.scala 189:26]
    .clock(mmioXbar_clock),
    .reset(mmioXbar_reset),
    .io_in_0_req_ready(mmioXbar_io_in_0_req_ready),
    .io_in_0_req_valid(mmioXbar_io_in_0_req_valid),
    .io_in_0_req_bits_addr(mmioXbar_io_in_0_req_bits_addr),
    .io_in_0_resp_valid(mmioXbar_io_in_0_resp_valid),
    .io_in_0_resp_bits_rdata(mmioXbar_io_in_0_resp_bits_rdata),
    .io_in_1_req_ready(mmioXbar_io_in_1_req_ready),
    .io_in_1_req_valid(mmioXbar_io_in_1_req_valid),
    .io_in_1_req_bits_addr(mmioXbar_io_in_1_req_bits_addr),
    .io_in_1_req_bits_size(mmioXbar_io_in_1_req_bits_size),
    .io_in_1_req_bits_cmd(mmioXbar_io_in_1_req_bits_cmd),
    .io_in_1_req_bits_wmask(mmioXbar_io_in_1_req_bits_wmask),
    .io_in_1_req_bits_wdata(mmioXbar_io_in_1_req_bits_wdata),
    .io_in_1_resp_valid(mmioXbar_io_in_1_resp_valid),
    .io_in_1_resp_bits_cmd(mmioXbar_io_in_1_resp_bits_cmd),
    .io_in_1_resp_bits_rdata(mmioXbar_io_in_1_resp_bits_rdata),
    .io_out_req_ready(mmioXbar_io_out_req_ready),
    .io_out_req_valid(mmioXbar_io_out_req_valid),
    .io_out_req_bits_addr(mmioXbar_io_out_req_bits_addr),
    .io_out_req_bits_size(mmioXbar_io_out_req_bits_size),
    .io_out_req_bits_cmd(mmioXbar_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(mmioXbar_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(mmioXbar_io_out_req_bits_wdata),
    .io_out_resp_ready(mmioXbar_io_out_resp_ready),
    .io_out_resp_valid(mmioXbar_io_out_resp_valid),
    .io_out_resp_bits_cmd(mmioXbar_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(mmioXbar_io_out_resp_bits_rdata)
  );
  SimpleBusCrossbarNto1_1 dmemXbar ( // @[src/main/scala/nutcore/NutCore.scala 190:26]
    .clock(dmemXbar_clock),
    .reset(dmemXbar_reset),
    .io_in_0_req_ready(dmemXbar_io_in_0_req_ready),
    .io_in_0_req_valid(dmemXbar_io_in_0_req_valid),
    .io_in_0_req_bits_addr(dmemXbar_io_in_0_req_bits_addr),
    .io_in_0_req_bits_size(dmemXbar_io_in_0_req_bits_size),
    .io_in_0_req_bits_cmd(dmemXbar_io_in_0_req_bits_cmd),
    .io_in_0_req_bits_wmask(dmemXbar_io_in_0_req_bits_wmask),
    .io_in_0_req_bits_wdata(dmemXbar_io_in_0_req_bits_wdata),
    .io_in_0_resp_valid(dmemXbar_io_in_0_resp_valid),
    .io_in_0_resp_bits_rdata(dmemXbar_io_in_0_resp_bits_rdata),
    .io_in_3_req_ready(dmemXbar_io_in_3_req_ready),
    .io_in_3_req_valid(dmemXbar_io_in_3_req_valid),
    .io_in_3_req_bits_addr(dmemXbar_io_in_3_req_bits_addr),
    .io_in_3_req_bits_size(dmemXbar_io_in_3_req_bits_size),
    .io_in_3_req_bits_cmd(dmemXbar_io_in_3_req_bits_cmd),
    .io_in_3_req_bits_wmask(dmemXbar_io_in_3_req_bits_wmask),
    .io_in_3_req_bits_wdata(dmemXbar_io_in_3_req_bits_wdata),
    .io_in_3_resp_ready(dmemXbar_io_in_3_resp_ready),
    .io_in_3_resp_valid(dmemXbar_io_in_3_resp_valid),
    .io_in_3_resp_bits_cmd(dmemXbar_io_in_3_resp_bits_cmd),
    .io_in_3_resp_bits_rdata(dmemXbar_io_in_3_resp_bits_rdata),
    .io_out_req_ready(dmemXbar_io_out_req_ready),
    .io_out_req_valid(dmemXbar_io_out_req_valid),
    .io_out_req_bits_addr(dmemXbar_io_out_req_bits_addr),
    .io_out_req_bits_size(dmemXbar_io_out_req_bits_size),
    .io_out_req_bits_cmd(dmemXbar_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(dmemXbar_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(dmemXbar_io_out_req_bits_wdata),
    .io_out_resp_ready(dmemXbar_io_out_resp_ready),
    .io_out_resp_valid(dmemXbar_io_out_resp_valid),
    .io_out_resp_bits_cmd(dmemXbar_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(dmemXbar_io_out_resp_bits_rdata)
  );
  EmbeddedTLB_fake itlb ( // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 438:13]
    .io_in_req_ready(itlb_io_in_req_ready),
    .io_in_req_valid(itlb_io_in_req_valid),
    .io_in_req_bits_addr(itlb_io_in_req_bits_addr),
    .io_in_req_bits_user(itlb_io_in_req_bits_user),
    .io_in_resp_ready(itlb_io_in_resp_ready),
    .io_in_resp_valid(itlb_io_in_resp_valid),
    .io_in_resp_bits_rdata(itlb_io_in_resp_bits_rdata),
    .io_in_resp_bits_user(itlb_io_in_resp_bits_user),
    .io_out_req_ready(itlb_io_out_req_ready),
    .io_out_req_valid(itlb_io_out_req_valid),
    .io_out_req_bits_addr(itlb_io_out_req_bits_addr),
    .io_out_req_bits_user(itlb_io_out_req_bits_user),
    .io_out_resp_ready(itlb_io_out_resp_ready),
    .io_out_resp_valid(itlb_io_out_resp_valid),
    .io_out_resp_bits_rdata(itlb_io_out_resp_bits_rdata),
    .io_out_resp_bits_user(itlb_io_out_resp_bits_user)
  );
  Cache_fake io_imem_cache ( // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
    .clock(io_imem_cache_clock),
    .reset(io_imem_cache_reset),
    .io_in_req_ready(io_imem_cache_io_in_req_ready),
    .io_in_req_valid(io_imem_cache_io_in_req_valid),
    .io_in_req_bits_addr(io_imem_cache_io_in_req_bits_addr),
    .io_in_req_bits_user(io_imem_cache_io_in_req_bits_user),
    .io_in_resp_ready(io_imem_cache_io_in_resp_ready),
    .io_in_resp_valid(io_imem_cache_io_in_resp_valid),
    .io_in_resp_bits_rdata(io_imem_cache_io_in_resp_bits_rdata),
    .io_in_resp_bits_user(io_imem_cache_io_in_resp_bits_user),
    .io_flush(io_imem_cache_io_flush),
    .io_out_mem_req_ready(io_imem_cache_io_out_mem_req_ready),
    .io_out_mem_req_valid(io_imem_cache_io_out_mem_req_valid),
    .io_out_mem_req_bits_addr(io_imem_cache_io_out_mem_req_bits_addr),
    .io_out_mem_resp_ready(io_imem_cache_io_out_mem_resp_ready),
    .io_out_mem_resp_valid(io_imem_cache_io_out_mem_resp_valid),
    .io_out_mem_resp_bits_rdata(io_imem_cache_io_out_mem_resp_bits_rdata),
    .io_mmio_req_ready(io_imem_cache_io_mmio_req_ready),
    .io_mmio_req_valid(io_imem_cache_io_mmio_req_valid),
    .io_mmio_req_bits_addr(io_imem_cache_io_mmio_req_bits_addr),
    .io_mmio_resp_ready(io_imem_cache_io_mmio_resp_ready),
    .io_mmio_resp_valid(io_imem_cache_io_mmio_resp_valid),
    .io_mmio_resp_bits_rdata(io_imem_cache_io_mmio_resp_bits_rdata)
  );
  EmbeddedTLB_fake_1 dtlb ( // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 438:13]
    .io_in_req_ready(dtlb_io_in_req_ready),
    .io_in_req_valid(dtlb_io_in_req_valid),
    .io_in_req_bits_addr(dtlb_io_in_req_bits_addr),
    .io_in_req_bits_size(dtlb_io_in_req_bits_size),
    .io_in_req_bits_cmd(dtlb_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(dtlb_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(dtlb_io_in_req_bits_wdata),
    .io_in_resp_valid(dtlb_io_in_resp_valid),
    .io_in_resp_bits_rdata(dtlb_io_in_resp_bits_rdata),
    .io_out_req_ready(dtlb_io_out_req_ready),
    .io_out_req_valid(dtlb_io_out_req_valid),
    .io_out_req_bits_addr(dtlb_io_out_req_bits_addr),
    .io_out_req_bits_size(dtlb_io_out_req_bits_size),
    .io_out_req_bits_cmd(dtlb_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(dtlb_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(dtlb_io_out_req_bits_wdata),
    .io_out_resp_valid(dtlb_io_out_resp_valid),
    .io_out_resp_bits_rdata(dtlb_io_out_resp_bits_rdata)
  );
  Cache_fake_1 io_dmem_cache ( // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
    .clock(io_dmem_cache_clock),
    .reset(io_dmem_cache_reset),
    .io_in_req_ready(io_dmem_cache_io_in_req_ready),
    .io_in_req_valid(io_dmem_cache_io_in_req_valid),
    .io_in_req_bits_addr(io_dmem_cache_io_in_req_bits_addr),
    .io_in_req_bits_size(io_dmem_cache_io_in_req_bits_size),
    .io_in_req_bits_cmd(io_dmem_cache_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(io_dmem_cache_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(io_dmem_cache_io_in_req_bits_wdata),
    .io_in_resp_ready(io_dmem_cache_io_in_resp_ready),
    .io_in_resp_valid(io_dmem_cache_io_in_resp_valid),
    .io_in_resp_bits_cmd(io_dmem_cache_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(io_dmem_cache_io_in_resp_bits_rdata),
    .io_out_mem_req_ready(io_dmem_cache_io_out_mem_req_ready),
    .io_out_mem_req_valid(io_dmem_cache_io_out_mem_req_valid),
    .io_out_mem_req_bits_addr(io_dmem_cache_io_out_mem_req_bits_addr),
    .io_out_mem_req_bits_size(io_dmem_cache_io_out_mem_req_bits_size),
    .io_out_mem_req_bits_cmd(io_dmem_cache_io_out_mem_req_bits_cmd),
    .io_out_mem_req_bits_wmask(io_dmem_cache_io_out_mem_req_bits_wmask),
    .io_out_mem_req_bits_wdata(io_dmem_cache_io_out_mem_req_bits_wdata),
    .io_out_mem_resp_ready(io_dmem_cache_io_out_mem_resp_ready),
    .io_out_mem_resp_valid(io_dmem_cache_io_out_mem_resp_valid),
    .io_out_mem_resp_bits_cmd(io_dmem_cache_io_out_mem_resp_bits_cmd),
    .io_out_mem_resp_bits_rdata(io_dmem_cache_io_out_mem_resp_bits_rdata),
    .io_mmio_req_ready(io_dmem_cache_io_mmio_req_ready),
    .io_mmio_req_valid(io_dmem_cache_io_mmio_req_valid),
    .io_mmio_req_bits_addr(io_dmem_cache_io_mmio_req_bits_addr),
    .io_mmio_req_bits_size(io_dmem_cache_io_mmio_req_bits_size),
    .io_mmio_req_bits_cmd(io_dmem_cache_io_mmio_req_bits_cmd),
    .io_mmio_req_bits_wmask(io_dmem_cache_io_mmio_req_bits_wmask),
    .io_mmio_req_bits_wdata(io_dmem_cache_io_mmio_req_bits_wdata),
    .io_mmio_resp_ready(io_dmem_cache_io_mmio_resp_ready),
    .io_mmio_resp_valid(io_dmem_cache_io_mmio_resp_valid),
    .io_mmio_resp_bits_cmd(io_dmem_cache_io_mmio_resp_bits_cmd),
    .io_mmio_resp_bits_rdata(io_dmem_cache_io_mmio_resp_bits_rdata)
  );
  assign io_imem_mem_req_valid = io_imem_cache_io_out_mem_req_valid; // @[src/main/scala/nutcore/NutCore.scala 194:13]
  assign io_imem_mem_req_bits_addr = io_imem_cache_io_out_mem_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 194:13]
  assign io_imem_mem_req_bits_size = 3'h3; // @[src/main/scala/nutcore/NutCore.scala 194:13]
  assign io_imem_mem_req_bits_cmd = 4'h0; // @[src/main/scala/nutcore/NutCore.scala 194:13]
  assign io_imem_mem_req_bits_wmask = 8'h0; // @[src/main/scala/nutcore/NutCore.scala 194:13]
  assign io_imem_mem_req_bits_wdata = 64'h0; // @[src/main/scala/nutcore/NutCore.scala 194:13]
  assign io_imem_mem_resp_ready = 1'h1; // @[src/main/scala/nutcore/NutCore.scala 194:13]
  assign io_imem_coh_req_ready = 1'h0; // @[src/main/scala/nutcore/NutCore.scala 194:13]
  assign io_imem_coh_resp_valid = 1'h0; // @[src/main/scala/nutcore/NutCore.scala 194:13]
  assign io_imem_coh_resp_bits_cmd = 4'h0; // @[src/main/scala/nutcore/NutCore.scala 194:13]
  assign io_imem_coh_resp_bits_rdata = 64'h0; // @[src/main/scala/nutcore/NutCore.scala 194:13]
  assign io_dmem_mem_req_valid = io_dmem_cache_io_out_mem_req_valid; // @[src/main/scala/nutcore/NutCore.scala 199:13]
  assign io_dmem_mem_req_bits_addr = io_dmem_cache_io_out_mem_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 199:13]
  assign io_dmem_mem_req_bits_size = io_dmem_cache_io_out_mem_req_bits_size; // @[src/main/scala/nutcore/NutCore.scala 199:13]
  assign io_dmem_mem_req_bits_cmd = io_dmem_cache_io_out_mem_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 199:13]
  assign io_dmem_mem_req_bits_wmask = io_dmem_cache_io_out_mem_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 199:13]
  assign io_dmem_mem_req_bits_wdata = io_dmem_cache_io_out_mem_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 199:13]
  assign io_dmem_mem_resp_ready = 1'h1; // @[src/main/scala/nutcore/NutCore.scala 199:13]
  assign io_dmem_coh_req_ready = 1'h0; // @[src/main/scala/nutcore/NutCore.scala 199:13]
  assign io_dmem_coh_resp_valid = 1'h0; // @[src/main/scala/nutcore/NutCore.scala 199:13]
  assign io_dmem_coh_resp_bits_cmd = 4'h0; // @[src/main/scala/nutcore/NutCore.scala 199:13]
  assign io_dmem_coh_resp_bits_rdata = 64'h0; // @[src/main/scala/nutcore/NutCore.scala 199:13]
  assign io_mmio_req_valid = mmioXbar_io_out_req_valid; // @[src/main/scala/nutcore/NutCore.scala 208:13]
  assign io_mmio_req_bits_addr = mmioXbar_io_out_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 208:13]
  assign io_mmio_req_bits_size = mmioXbar_io_out_req_bits_size; // @[src/main/scala/nutcore/NutCore.scala 208:13]
  assign io_mmio_req_bits_cmd = mmioXbar_io_out_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 208:13]
  assign io_mmio_req_bits_wmask = mmioXbar_io_out_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 208:13]
  assign io_mmio_req_bits_wdata = mmioXbar_io_out_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 208:13]
  assign io_mmio_resp_ready = 1'h1; // @[src/main/scala/nutcore/NutCore.scala 208:13]
  assign io_frontend_req_ready = dmemXbar_io_in_3_req_ready; // @[src/main/scala/nutcore/NutCore.scala 206:23]
  assign io_frontend_resp_valid = dmemXbar_io_in_3_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 206:23]
  assign io_frontend_resp_bits_cmd = dmemXbar_io_in_3_resp_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 206:23]
  assign io_frontend_resp_bits_rdata = dmemXbar_io_in_3_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 206:23]
  assign rvfi_valid = backend_io_in_valid;
  assign rvfi_order = backend_rvfi_order;
  assign rvfi_insn = backend_io_in_bits_decode_cf_instr;
  assign rvfi_trap = backend_REG_0;
  assign rvfi_halt = 1'h0; // @[src/main/scala/nutcore/NutCore.scala 218:17]
  assign rvfi_intr = 1'h0; // @[src/main/scala/nutcore/NutCore.scala 219:17]
  assign rvfi_mode = 2'h3; // @[src/main/scala/nutcore/NutCore.scala 220:17]
  assign rvfi_ixl = 2'h1; // @[src/main/scala/nutcore/NutCore.scala 221:17]
  assign rvfi_rs1_addr = backend_io_in_bits_decode_ctrl_rfSrc1;
  assign rvfi_rs2_addr = backend_io_in_bits_decode_ctrl_rfSrc2;
  assign rvfi_rs1_rdata = backend_io_in_bits_decode_data_src1;
  assign rvfi_rs2_rdata = backend_io_in_bits_decode_data_src2;
  assign rvfi_rd_addr = backend_io_wb_rfDest;
  assign rvfi_rd_wdata = backend__T_142;
  assign rvfi_pc_rdata = backend__T_145;
  assign rvfi_pc_wdata = backend__T_151;
  assign rvfi_mem_addr = {_rvfi_mem_addr_T_4,_rvfi_mem_addr_T_2}; // @[src/main/scala/utils/BitUtils.scala 40:41]
  assign rvfi_mem_rmask = backend_io_in_bits_mem_rvfi_rmask;
  assign rvfi_mem_wmask = backend_io_in_bits_mem_rvfi_wmask;
  assign rvfi_mem_rdata = backend_io_in_bits_mem_rvfi_rdata;
  assign rvfi_mem_wdata = backend_io_in_bits_mem_rvfi_wdata;
  assign frontend_clock = clock;
  assign frontend_reset = reset;
  assign frontend_io_imem_req_ready = itlb_io_in_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 440:15]
  assign frontend_io_imem_resp_valid = itlb_io_in_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 440:15]
  assign frontend_io_imem_resp_bits_rdata = itlb_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 440:15]
  assign frontend_io_imem_resp_bits_user = itlb_io_in_resp_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 440:15]
  assign frontend_io_out_0_ready = ringBufferAllowin | ~frontend_io_out_0_valid; // @[src/main/scala/utils/PipelineVector.scala 50:36]
  assign frontend_io_redirect_target = backend_io_redirect_target; // @[src/main/scala/nutcore/NutCore.scala 202:26]
  assign frontend_io_redirect_valid = backend_io_redirect_valid; // @[src/main/scala/nutcore/NutCore.scala 202:26]
  assign frontend_flushICache = backend_flushICache;
  assign frontend_REG_valid = backend_REG_valid;
  assign frontend_REG_pc = backend_REG_pc;
  assign frontend_REG_isMissPredict = backend_REG_isMissPredict;
  assign frontend_REG_actualTarget = backend_REG_actualTarget;
  assign frontend_REG_actualTaken = backend_REG_actualTaken;
  assign frontend_REG_fuOpType = backend_REG_fuOpType;
  assign frontend_REG_btbType = backend_REG_btbType;
  assign frontend_REG_isRVC = backend_REG_isRVC;
  assign frontend_intrVec = backend_intrVec;
  assign frontend_flushTLB = backend_flushTLB;
  assign backend_clock = clock;
  assign backend_reset = reset;
  assign backend_io_in_0_valid = ringBufferHead != ringBufferTail; // @[src/main/scala/utils/PipelineVector.scala 56:34]
  assign backend_io_in_0_bits_cf_instr = 2'h3 == ringBufferTail ? dataBuffer_3_cf_instr : _GEN_1319; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_pc = 2'h3 == ringBufferTail ? dataBuffer_3_cf_pc : _GEN_1315; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_pnpc = 2'h3 == ringBufferTail ? dataBuffer_3_cf_pnpc : _GEN_1311; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_exceptionVec_1 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_exceptionVec_1 : _GEN_1239; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_exceptionVec_2 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_exceptionVec_2 : _GEN_1243; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_0 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_intrVec_0 : _GEN_1187; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_1 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_intrVec_1 : _GEN_1191; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_2 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_intrVec_2 : _GEN_1195; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_3 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_intrVec_3 : _GEN_1199; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_4 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_intrVec_4 : _GEN_1203; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_5 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_intrVec_5 : _GEN_1207; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_6 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_intrVec_6 : _GEN_1211; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_7 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_intrVec_7 : _GEN_1215; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_8 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_intrVec_8 : _GEN_1219; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_9 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_intrVec_9 : _GEN_1223; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_10 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_intrVec_10 : _GEN_1227; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_11 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_intrVec_11 : _GEN_1231; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_brIdx = 2'h3 == ringBufferTail ? dataBuffer_3_cf_brIdx : _GEN_1183; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_src1Type = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_src1Type : _GEN_1163; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_src2Type = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_src2Type : _GEN_1159; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_fuType = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_fuType : _GEN_1155; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_fuOpType = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_fuOpType : _GEN_1151; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_rfSrc1 = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_rfSrc1 : _GEN_1147; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_rfSrc2 = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_rfSrc2 : _GEN_1143; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_rfWen = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_rfWen : _GEN_1139; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_rfDest = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_rfDest : _GEN_1135; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_data_imm = 2'h3 == ringBufferTail ? dataBuffer_3_data_imm : _GEN_1103; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_flush = frontend_io_flushVec[3:2]; // @[src/main/scala/nutcore/NutCore.scala 203:45]
  assign backend_io_dmem_req_ready = dtlb_io_in_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 440:15]
  assign backend_io_dmem_resp_valid = dtlb_io_in_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 440:15]
  assign backend_io_dmem_resp_bits_rdata = dtlb_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 440:15]
  assign mmioXbar_clock = clock;
  assign mmioXbar_reset = reset;
  assign mmioXbar_io_in_0_req_valid = io_imem_cache_io_mmio_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign mmioXbar_io_in_0_req_bits_addr = io_imem_cache_io_mmio_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign mmioXbar_io_in_1_req_valid = io_dmem_cache_io_mmio_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign mmioXbar_io_in_1_req_bits_addr = io_dmem_cache_io_mmio_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign mmioXbar_io_in_1_req_bits_size = io_dmem_cache_io_mmio_req_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign mmioXbar_io_in_1_req_bits_cmd = io_dmem_cache_io_mmio_req_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign mmioXbar_io_in_1_req_bits_wmask = io_dmem_cache_io_mmio_req_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign mmioXbar_io_in_1_req_bits_wdata = io_dmem_cache_io_mmio_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign mmioXbar_io_out_req_ready = io_mmio_req_ready; // @[src/main/scala/nutcore/NutCore.scala 208:13]
  assign mmioXbar_io_out_resp_valid = io_mmio_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 208:13]
  assign mmioXbar_io_out_resp_bits_cmd = io_mmio_resp_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 208:13]
  assign mmioXbar_io_out_resp_bits_rdata = io_mmio_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 208:13]
  assign dmemXbar_clock = clock;
  assign dmemXbar_reset = reset;
  assign dmemXbar_io_in_0_req_valid = dtlb_io_out_req_valid; // @[src/main/scala/nutcore/NutCore.scala 198:23]
  assign dmemXbar_io_in_0_req_bits_addr = dtlb_io_out_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 198:23]
  assign dmemXbar_io_in_0_req_bits_size = dtlb_io_out_req_bits_size; // @[src/main/scala/nutcore/NutCore.scala 198:23]
  assign dmemXbar_io_in_0_req_bits_cmd = dtlb_io_out_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 198:23]
  assign dmemXbar_io_in_0_req_bits_wmask = dtlb_io_out_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 198:23]
  assign dmemXbar_io_in_0_req_bits_wdata = dtlb_io_out_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 198:23]
  assign dmemXbar_io_in_3_req_valid = io_frontend_req_valid; // @[src/main/scala/nutcore/NutCore.scala 206:23]
  assign dmemXbar_io_in_3_req_bits_addr = io_frontend_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 206:23]
  assign dmemXbar_io_in_3_req_bits_size = io_frontend_req_bits_size; // @[src/main/scala/nutcore/NutCore.scala 206:23]
  assign dmemXbar_io_in_3_req_bits_cmd = io_frontend_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 206:23]
  assign dmemXbar_io_in_3_req_bits_wmask = io_frontend_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 206:23]
  assign dmemXbar_io_in_3_req_bits_wdata = io_frontend_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 206:23]
  assign dmemXbar_io_in_3_resp_ready = io_frontend_resp_ready; // @[src/main/scala/nutcore/NutCore.scala 206:23]
  assign dmemXbar_io_out_req_ready = io_dmem_cache_io_in_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign dmemXbar_io_out_resp_valid = io_dmem_cache_io_in_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign dmemXbar_io_out_resp_bits_cmd = io_dmem_cache_io_in_resp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign dmemXbar_io_out_resp_bits_rdata = io_dmem_cache_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign itlb_io_in_req_valid = frontend_io_imem_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 440:15]
  assign itlb_io_in_req_bits_addr = frontend_io_imem_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 440:15]
  assign itlb_io_in_req_bits_user = frontend_io_imem_req_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 440:15]
  assign itlb_io_in_resp_ready = frontend_io_imem_resp_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 440:15]
  assign itlb_io_out_req_ready = io_imem_cache_io_in_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign itlb_io_out_resp_valid = io_imem_cache_io_in_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign itlb_io_out_resp_bits_rdata = io_imem_cache_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign itlb_io_out_resp_bits_user = io_imem_cache_io_in_resp_bits_user; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign io_imem_cache_clock = clock;
  assign io_imem_cache_reset = reset;
  assign io_imem_cache_io_in_req_valid = itlb_io_out_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign io_imem_cache_io_in_req_bits_addr = itlb_io_out_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign io_imem_cache_io_in_req_bits_user = itlb_io_out_req_bits_user; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign io_imem_cache_io_in_resp_ready = itlb_io_out_resp_ready; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign io_imem_cache_io_flush = frontend_io_flushVec[0] ? 2'h3 : 2'h0; // @[src/main/scala/nutcore/NutCore.scala 194:83]
  assign io_imem_cache_io_out_mem_req_ready = io_imem_mem_req_ready; // @[src/main/scala/nutcore/NutCore.scala 194:13]
  assign io_imem_cache_io_out_mem_resp_valid = io_imem_mem_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 194:13]
  assign io_imem_cache_io_out_mem_resp_bits_rdata = io_imem_mem_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 194:13]
  assign io_imem_cache_io_mmio_req_ready = mmioXbar_io_in_0_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign io_imem_cache_io_mmio_resp_valid = mmioXbar_io_in_0_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign io_imem_cache_io_mmio_resp_bits_rdata = mmioXbar_io_in_0_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign dtlb_io_in_req_valid = backend_io_dmem_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 440:15]
  assign dtlb_io_in_req_bits_addr = backend_io_dmem_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 440:15]
  assign dtlb_io_in_req_bits_size = backend_io_dmem_req_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 440:15]
  assign dtlb_io_in_req_bits_cmd = backend_io_dmem_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 440:15]
  assign dtlb_io_in_req_bits_wmask = backend_io_dmem_req_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 440:15]
  assign dtlb_io_in_req_bits_wdata = backend_io_dmem_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 440:15]
  assign dtlb_io_out_req_ready = dmemXbar_io_in_0_req_ready; // @[src/main/scala/nutcore/NutCore.scala 198:23]
  assign dtlb_io_out_resp_valid = dmemXbar_io_in_0_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 198:23]
  assign dtlb_io_out_resp_bits_rdata = dmemXbar_io_in_0_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 198:23]
  assign io_dmem_cache_clock = clock;
  assign io_dmem_cache_reset = reset;
  assign io_dmem_cache_io_in_req_valid = dmemXbar_io_out_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign io_dmem_cache_io_in_req_bits_addr = dmemXbar_io_out_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign io_dmem_cache_io_in_req_bits_size = dmemXbar_io_out_req_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign io_dmem_cache_io_in_req_bits_cmd = dmemXbar_io_out_req_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign io_dmem_cache_io_in_req_bits_wmask = dmemXbar_io_out_req_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign io_dmem_cache_io_in_req_bits_wdata = dmemXbar_io_out_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign io_dmem_cache_io_in_resp_ready = dmemXbar_io_out_resp_ready; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign io_dmem_cache_io_out_mem_req_ready = io_dmem_mem_req_ready; // @[src/main/scala/nutcore/NutCore.scala 199:13]
  assign io_dmem_cache_io_out_mem_resp_valid = io_dmem_mem_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 199:13]
  assign io_dmem_cache_io_out_mem_resp_bits_cmd = io_dmem_mem_resp_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 199:13]
  assign io_dmem_cache_io_out_mem_resp_bits_rdata = io_dmem_mem_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 199:13]
  assign io_dmem_cache_io_mmio_req_ready = mmioXbar_io_in_1_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign io_dmem_cache_io_mmio_resp_valid = mmioXbar_io_in_1_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign io_dmem_cache_io_mmio_resp_bits_cmd = mmioXbar_io_in_1_resp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign io_dmem_cache_io_mmio_resp_bits_rdata = mmioXbar_io_in_1_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_instr <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_instr <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_instr <= _GEN_220;
        end
      end else begin
        dataBuffer_0_cf_instr <= _GEN_220;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_pc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_pc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_pc <= _GEN_224;
        end
      end else begin
        dataBuffer_0_cf_pc <= _GEN_224;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_pnpc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_pnpc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_pnpc <= _GEN_228;
        end
      end else begin
        dataBuffer_0_cf_pnpc <= _GEN_228;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_exceptionVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_exceptionVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_exceptionVec_1 <= _GEN_248;
        end
      end else begin
        dataBuffer_0_cf_exceptionVec_1 <= _GEN_248;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_exceptionVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_exceptionVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_exceptionVec_2 <= _GEN_252;
        end
      end else begin
        dataBuffer_0_cf_exceptionVec_2 <= _GEN_252;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_intrVec_0 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_intrVec_0 <= frontend_io_out_1_bits_cf_intrVec_0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_intrVec_0 <= _GEN_308;
        end
      end else begin
        dataBuffer_0_cf_intrVec_0 <= _GEN_308;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_intrVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_intrVec_1 <= frontend_io_out_1_bits_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_intrVec_1 <= _GEN_312;
        end
      end else begin
        dataBuffer_0_cf_intrVec_1 <= _GEN_312;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_intrVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_intrVec_2 <= frontend_io_out_1_bits_cf_intrVec_2; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_intrVec_2 <= _GEN_316;
        end
      end else begin
        dataBuffer_0_cf_intrVec_2 <= _GEN_316;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_intrVec_3 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_intrVec_3 <= frontend_io_out_1_bits_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_intrVec_3 <= _GEN_320;
        end
      end else begin
        dataBuffer_0_cf_intrVec_3 <= _GEN_320;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_intrVec_4 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_intrVec_4 <= frontend_io_out_1_bits_cf_intrVec_4; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_intrVec_4 <= _GEN_324;
        end
      end else begin
        dataBuffer_0_cf_intrVec_4 <= _GEN_324;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_intrVec_5 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_intrVec_5 <= frontend_io_out_1_bits_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_intrVec_5 <= _GEN_328;
        end
      end else begin
        dataBuffer_0_cf_intrVec_5 <= _GEN_328;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_intrVec_6 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_intrVec_6 <= frontend_io_out_1_bits_cf_intrVec_6; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_intrVec_6 <= _GEN_332;
        end
      end else begin
        dataBuffer_0_cf_intrVec_6 <= _GEN_332;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_intrVec_7 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_intrVec_7 <= frontend_io_out_1_bits_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_intrVec_7 <= _GEN_336;
        end
      end else begin
        dataBuffer_0_cf_intrVec_7 <= _GEN_336;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_intrVec_8 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_intrVec_8 <= frontend_io_out_1_bits_cf_intrVec_8; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_intrVec_8 <= _GEN_340;
        end
      end else begin
        dataBuffer_0_cf_intrVec_8 <= _GEN_340;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_intrVec_9 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_intrVec_9 <= frontend_io_out_1_bits_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_intrVec_9 <= _GEN_344;
        end
      end else begin
        dataBuffer_0_cf_intrVec_9 <= _GEN_344;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_intrVec_10 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_intrVec_10 <= frontend_io_out_1_bits_cf_intrVec_10; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_intrVec_10 <= _GEN_348;
        end
      end else begin
        dataBuffer_0_cf_intrVec_10 <= _GEN_348;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_intrVec_11 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_intrVec_11 <= frontend_io_out_1_bits_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_intrVec_11 <= _GEN_352;
        end
      end else begin
        dataBuffer_0_cf_intrVec_11 <= _GEN_352;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_brIdx <= 4'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_brIdx <= 4'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_brIdx <= _GEN_356;
        end
      end else begin
        dataBuffer_0_cf_brIdx <= _GEN_356;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_src1Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        dataBuffer_0_ctrl_src1Type <= 2'h0 == _T_7 | _GEN_376;
      end else if (enqueueFire_0) begin // @[src/main/scala/utils/PipelineVector.scala 45:29]
        dataBuffer_0_ctrl_src1Type <= _GEN_156;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_src2Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        dataBuffer_0_ctrl_src2Type <= 2'h0 == _T_7 | _GEN_380;
      end else if (enqueueFire_0) begin // @[src/main/scala/utils/PipelineVector.scala 45:29]
        dataBuffer_0_ctrl_src2Type <= _GEN_160;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_fuType <= 3'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_ctrl_fuType <= 3'h3; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_ctrl_fuType <= _GEN_384;
        end
      end else begin
        dataBuffer_0_ctrl_fuType <= _GEN_384;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_fuOpType <= 7'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_ctrl_fuOpType <= 7'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_ctrl_fuOpType <= _GEN_388;
        end
      end else begin
        dataBuffer_0_ctrl_fuOpType <= _GEN_388;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_rfSrc1 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_ctrl_rfSrc1 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_ctrl_rfSrc1 <= _GEN_392;
        end
      end else begin
        dataBuffer_0_ctrl_rfSrc1 <= _GEN_392;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_rfSrc2 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_ctrl_rfSrc2 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_ctrl_rfSrc2 <= _GEN_396;
        end
      end else begin
        dataBuffer_0_ctrl_rfSrc2 <= _GEN_396;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_rfWen <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_ctrl_rfWen <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_ctrl_rfWen <= _GEN_400;
        end
      end else begin
        dataBuffer_0_ctrl_rfWen <= _GEN_400;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_rfDest <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_ctrl_rfDest <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_ctrl_rfDest <= _GEN_404;
        end
      end else begin
        dataBuffer_0_ctrl_rfDest <= _GEN_404;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_data_imm <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_data_imm <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_data_imm <= _GEN_436;
        end
      end else begin
        dataBuffer_0_data_imm <= _GEN_436;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_instr <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_instr <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_instr <= _GEN_221;
        end
      end else begin
        dataBuffer_1_cf_instr <= _GEN_221;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_pc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_pc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_pc <= _GEN_225;
        end
      end else begin
        dataBuffer_1_cf_pc <= _GEN_225;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_pnpc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_pnpc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_pnpc <= _GEN_229;
        end
      end else begin
        dataBuffer_1_cf_pnpc <= _GEN_229;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_exceptionVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_exceptionVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_exceptionVec_1 <= _GEN_249;
        end
      end else begin
        dataBuffer_1_cf_exceptionVec_1 <= _GEN_249;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_exceptionVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_exceptionVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_exceptionVec_2 <= _GEN_253;
        end
      end else begin
        dataBuffer_1_cf_exceptionVec_2 <= _GEN_253;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_intrVec_0 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_intrVec_0 <= frontend_io_out_1_bits_cf_intrVec_0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_intrVec_0 <= _GEN_309;
        end
      end else begin
        dataBuffer_1_cf_intrVec_0 <= _GEN_309;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_intrVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_intrVec_1 <= frontend_io_out_1_bits_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_intrVec_1 <= _GEN_313;
        end
      end else begin
        dataBuffer_1_cf_intrVec_1 <= _GEN_313;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_intrVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_intrVec_2 <= frontend_io_out_1_bits_cf_intrVec_2; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_intrVec_2 <= _GEN_317;
        end
      end else begin
        dataBuffer_1_cf_intrVec_2 <= _GEN_317;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_intrVec_3 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_intrVec_3 <= frontend_io_out_1_bits_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_intrVec_3 <= _GEN_321;
        end
      end else begin
        dataBuffer_1_cf_intrVec_3 <= _GEN_321;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_intrVec_4 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_intrVec_4 <= frontend_io_out_1_bits_cf_intrVec_4; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_intrVec_4 <= _GEN_325;
        end
      end else begin
        dataBuffer_1_cf_intrVec_4 <= _GEN_325;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_intrVec_5 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_intrVec_5 <= frontend_io_out_1_bits_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_intrVec_5 <= _GEN_329;
        end
      end else begin
        dataBuffer_1_cf_intrVec_5 <= _GEN_329;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_intrVec_6 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_intrVec_6 <= frontend_io_out_1_bits_cf_intrVec_6; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_intrVec_6 <= _GEN_333;
        end
      end else begin
        dataBuffer_1_cf_intrVec_6 <= _GEN_333;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_intrVec_7 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_intrVec_7 <= frontend_io_out_1_bits_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_intrVec_7 <= _GEN_337;
        end
      end else begin
        dataBuffer_1_cf_intrVec_7 <= _GEN_337;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_intrVec_8 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_intrVec_8 <= frontend_io_out_1_bits_cf_intrVec_8; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_intrVec_8 <= _GEN_341;
        end
      end else begin
        dataBuffer_1_cf_intrVec_8 <= _GEN_341;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_intrVec_9 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_intrVec_9 <= frontend_io_out_1_bits_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_intrVec_9 <= _GEN_345;
        end
      end else begin
        dataBuffer_1_cf_intrVec_9 <= _GEN_345;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_intrVec_10 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_intrVec_10 <= frontend_io_out_1_bits_cf_intrVec_10; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_intrVec_10 <= _GEN_349;
        end
      end else begin
        dataBuffer_1_cf_intrVec_10 <= _GEN_349;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_intrVec_11 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_intrVec_11 <= frontend_io_out_1_bits_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_intrVec_11 <= _GEN_353;
        end
      end else begin
        dataBuffer_1_cf_intrVec_11 <= _GEN_353;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_brIdx <= 4'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_brIdx <= 4'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_brIdx <= _GEN_357;
        end
      end else begin
        dataBuffer_1_cf_brIdx <= _GEN_357;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_src1Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        dataBuffer_1_ctrl_src1Type <= 2'h1 == _T_7 | _GEN_377;
      end else if (enqueueFire_0) begin // @[src/main/scala/utils/PipelineVector.scala 45:29]
        dataBuffer_1_ctrl_src1Type <= _GEN_157;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_src2Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        dataBuffer_1_ctrl_src2Type <= 2'h1 == _T_7 | _GEN_381;
      end else if (enqueueFire_0) begin // @[src/main/scala/utils/PipelineVector.scala 45:29]
        dataBuffer_1_ctrl_src2Type <= _GEN_161;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_fuType <= 3'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_ctrl_fuType <= 3'h3; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_ctrl_fuType <= _GEN_385;
        end
      end else begin
        dataBuffer_1_ctrl_fuType <= _GEN_385;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_fuOpType <= 7'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_ctrl_fuOpType <= 7'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_ctrl_fuOpType <= _GEN_389;
        end
      end else begin
        dataBuffer_1_ctrl_fuOpType <= _GEN_389;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_rfSrc1 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_ctrl_rfSrc1 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_ctrl_rfSrc1 <= _GEN_393;
        end
      end else begin
        dataBuffer_1_ctrl_rfSrc1 <= _GEN_393;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_rfSrc2 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_ctrl_rfSrc2 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_ctrl_rfSrc2 <= _GEN_397;
        end
      end else begin
        dataBuffer_1_ctrl_rfSrc2 <= _GEN_397;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_rfWen <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_ctrl_rfWen <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_ctrl_rfWen <= _GEN_401;
        end
      end else begin
        dataBuffer_1_ctrl_rfWen <= _GEN_401;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_rfDest <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_ctrl_rfDest <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_ctrl_rfDest <= _GEN_405;
        end
      end else begin
        dataBuffer_1_ctrl_rfDest <= _GEN_405;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_data_imm <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_data_imm <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_data_imm <= _GEN_437;
        end
      end else begin
        dataBuffer_1_data_imm <= _GEN_437;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_instr <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_instr <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_instr <= _GEN_222;
        end
      end else begin
        dataBuffer_2_cf_instr <= _GEN_222;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_pc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_pc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_pc <= _GEN_226;
        end
      end else begin
        dataBuffer_2_cf_pc <= _GEN_226;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_pnpc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_pnpc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_pnpc <= _GEN_230;
        end
      end else begin
        dataBuffer_2_cf_pnpc <= _GEN_230;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_exceptionVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_exceptionVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_exceptionVec_1 <= _GEN_250;
        end
      end else begin
        dataBuffer_2_cf_exceptionVec_1 <= _GEN_250;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_exceptionVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_exceptionVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_exceptionVec_2 <= _GEN_254;
        end
      end else begin
        dataBuffer_2_cf_exceptionVec_2 <= _GEN_254;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_intrVec_0 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_intrVec_0 <= frontend_io_out_1_bits_cf_intrVec_0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_intrVec_0 <= _GEN_310;
        end
      end else begin
        dataBuffer_2_cf_intrVec_0 <= _GEN_310;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_intrVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_intrVec_1 <= frontend_io_out_1_bits_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_intrVec_1 <= _GEN_314;
        end
      end else begin
        dataBuffer_2_cf_intrVec_1 <= _GEN_314;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_intrVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_intrVec_2 <= frontend_io_out_1_bits_cf_intrVec_2; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_intrVec_2 <= _GEN_318;
        end
      end else begin
        dataBuffer_2_cf_intrVec_2 <= _GEN_318;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_intrVec_3 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_intrVec_3 <= frontend_io_out_1_bits_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_intrVec_3 <= _GEN_322;
        end
      end else begin
        dataBuffer_2_cf_intrVec_3 <= _GEN_322;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_intrVec_4 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_intrVec_4 <= frontend_io_out_1_bits_cf_intrVec_4; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_intrVec_4 <= _GEN_326;
        end
      end else begin
        dataBuffer_2_cf_intrVec_4 <= _GEN_326;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_intrVec_5 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_intrVec_5 <= frontend_io_out_1_bits_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_intrVec_5 <= _GEN_330;
        end
      end else begin
        dataBuffer_2_cf_intrVec_5 <= _GEN_330;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_intrVec_6 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_intrVec_6 <= frontend_io_out_1_bits_cf_intrVec_6; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_intrVec_6 <= _GEN_334;
        end
      end else begin
        dataBuffer_2_cf_intrVec_6 <= _GEN_334;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_intrVec_7 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_intrVec_7 <= frontend_io_out_1_bits_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_intrVec_7 <= _GEN_338;
        end
      end else begin
        dataBuffer_2_cf_intrVec_7 <= _GEN_338;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_intrVec_8 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_intrVec_8 <= frontend_io_out_1_bits_cf_intrVec_8; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_intrVec_8 <= _GEN_342;
        end
      end else begin
        dataBuffer_2_cf_intrVec_8 <= _GEN_342;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_intrVec_9 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_intrVec_9 <= frontend_io_out_1_bits_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_intrVec_9 <= _GEN_346;
        end
      end else begin
        dataBuffer_2_cf_intrVec_9 <= _GEN_346;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_intrVec_10 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_intrVec_10 <= frontend_io_out_1_bits_cf_intrVec_10; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_intrVec_10 <= _GEN_350;
        end
      end else begin
        dataBuffer_2_cf_intrVec_10 <= _GEN_350;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_intrVec_11 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_intrVec_11 <= frontend_io_out_1_bits_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_intrVec_11 <= _GEN_354;
        end
      end else begin
        dataBuffer_2_cf_intrVec_11 <= _GEN_354;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_brIdx <= 4'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_brIdx <= 4'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_brIdx <= _GEN_358;
        end
      end else begin
        dataBuffer_2_cf_brIdx <= _GEN_358;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_src1Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        dataBuffer_2_ctrl_src1Type <= 2'h2 == _T_7 | _GEN_378;
      end else if (enqueueFire_0) begin // @[src/main/scala/utils/PipelineVector.scala 45:29]
        dataBuffer_2_ctrl_src1Type <= _GEN_158;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_src2Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        dataBuffer_2_ctrl_src2Type <= 2'h2 == _T_7 | _GEN_382;
      end else if (enqueueFire_0) begin // @[src/main/scala/utils/PipelineVector.scala 45:29]
        dataBuffer_2_ctrl_src2Type <= _GEN_162;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_fuType <= 3'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_ctrl_fuType <= 3'h3; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_ctrl_fuType <= _GEN_386;
        end
      end else begin
        dataBuffer_2_ctrl_fuType <= _GEN_386;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_fuOpType <= 7'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_ctrl_fuOpType <= 7'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_ctrl_fuOpType <= _GEN_390;
        end
      end else begin
        dataBuffer_2_ctrl_fuOpType <= _GEN_390;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_rfSrc1 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_ctrl_rfSrc1 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_ctrl_rfSrc1 <= _GEN_394;
        end
      end else begin
        dataBuffer_2_ctrl_rfSrc1 <= _GEN_394;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_rfSrc2 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_ctrl_rfSrc2 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_ctrl_rfSrc2 <= _GEN_398;
        end
      end else begin
        dataBuffer_2_ctrl_rfSrc2 <= _GEN_398;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_rfWen <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_ctrl_rfWen <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_ctrl_rfWen <= _GEN_402;
        end
      end else begin
        dataBuffer_2_ctrl_rfWen <= _GEN_402;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_rfDest <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_ctrl_rfDest <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_ctrl_rfDest <= _GEN_406;
        end
      end else begin
        dataBuffer_2_ctrl_rfDest <= _GEN_406;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_data_imm <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_data_imm <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_data_imm <= _GEN_438;
        end
      end else begin
        dataBuffer_2_data_imm <= _GEN_438;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_instr <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_instr <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_instr <= _GEN_223;
        end
      end else begin
        dataBuffer_3_cf_instr <= _GEN_223;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_pc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_pc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_pc <= _GEN_227;
        end
      end else begin
        dataBuffer_3_cf_pc <= _GEN_227;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_pnpc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_pnpc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_pnpc <= _GEN_231;
        end
      end else begin
        dataBuffer_3_cf_pnpc <= _GEN_231;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_exceptionVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_exceptionVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_exceptionVec_1 <= _GEN_251;
        end
      end else begin
        dataBuffer_3_cf_exceptionVec_1 <= _GEN_251;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_exceptionVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_exceptionVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_exceptionVec_2 <= _GEN_255;
        end
      end else begin
        dataBuffer_3_cf_exceptionVec_2 <= _GEN_255;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_intrVec_0 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_intrVec_0 <= frontend_io_out_1_bits_cf_intrVec_0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_intrVec_0 <= _GEN_311;
        end
      end else begin
        dataBuffer_3_cf_intrVec_0 <= _GEN_311;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_intrVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_intrVec_1 <= frontend_io_out_1_bits_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_intrVec_1 <= _GEN_315;
        end
      end else begin
        dataBuffer_3_cf_intrVec_1 <= _GEN_315;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_intrVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_intrVec_2 <= frontend_io_out_1_bits_cf_intrVec_2; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_intrVec_2 <= _GEN_319;
        end
      end else begin
        dataBuffer_3_cf_intrVec_2 <= _GEN_319;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_intrVec_3 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_intrVec_3 <= frontend_io_out_1_bits_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_intrVec_3 <= _GEN_323;
        end
      end else begin
        dataBuffer_3_cf_intrVec_3 <= _GEN_323;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_intrVec_4 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_intrVec_4 <= frontend_io_out_1_bits_cf_intrVec_4; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_intrVec_4 <= _GEN_327;
        end
      end else begin
        dataBuffer_3_cf_intrVec_4 <= _GEN_327;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_intrVec_5 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_intrVec_5 <= frontend_io_out_1_bits_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_intrVec_5 <= _GEN_331;
        end
      end else begin
        dataBuffer_3_cf_intrVec_5 <= _GEN_331;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_intrVec_6 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_intrVec_6 <= frontend_io_out_1_bits_cf_intrVec_6; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_intrVec_6 <= _GEN_335;
        end
      end else begin
        dataBuffer_3_cf_intrVec_6 <= _GEN_335;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_intrVec_7 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_intrVec_7 <= frontend_io_out_1_bits_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_intrVec_7 <= _GEN_339;
        end
      end else begin
        dataBuffer_3_cf_intrVec_7 <= _GEN_339;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_intrVec_8 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_intrVec_8 <= frontend_io_out_1_bits_cf_intrVec_8; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_intrVec_8 <= _GEN_343;
        end
      end else begin
        dataBuffer_3_cf_intrVec_8 <= _GEN_343;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_intrVec_9 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_intrVec_9 <= frontend_io_out_1_bits_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_intrVec_9 <= _GEN_347;
        end
      end else begin
        dataBuffer_3_cf_intrVec_9 <= _GEN_347;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_intrVec_10 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_intrVec_10 <= frontend_io_out_1_bits_cf_intrVec_10; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_intrVec_10 <= _GEN_351;
        end
      end else begin
        dataBuffer_3_cf_intrVec_10 <= _GEN_351;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_intrVec_11 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_intrVec_11 <= frontend_io_out_1_bits_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_intrVec_11 <= _GEN_355;
        end
      end else begin
        dataBuffer_3_cf_intrVec_11 <= _GEN_355;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_brIdx <= 4'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_brIdx <= 4'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_brIdx <= _GEN_359;
        end
      end else begin
        dataBuffer_3_cf_brIdx <= _GEN_359;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_src1Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        dataBuffer_3_ctrl_src1Type <= 2'h3 == _T_7 | _GEN_379;
      end else if (enqueueFire_0) begin // @[src/main/scala/utils/PipelineVector.scala 45:29]
        dataBuffer_3_ctrl_src1Type <= _GEN_159;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_src2Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        dataBuffer_3_ctrl_src2Type <= 2'h3 == _T_7 | _GEN_383;
      end else if (enqueueFire_0) begin // @[src/main/scala/utils/PipelineVector.scala 45:29]
        dataBuffer_3_ctrl_src2Type <= _GEN_163;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_fuType <= 3'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_ctrl_fuType <= 3'h3; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_ctrl_fuType <= _GEN_387;
        end
      end else begin
        dataBuffer_3_ctrl_fuType <= _GEN_387;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_fuOpType <= 7'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_ctrl_fuOpType <= 7'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_ctrl_fuOpType <= _GEN_391;
        end
      end else begin
        dataBuffer_3_ctrl_fuOpType <= _GEN_391;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_rfSrc1 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_ctrl_rfSrc1 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_ctrl_rfSrc1 <= _GEN_395;
        end
      end else begin
        dataBuffer_3_ctrl_rfSrc1 <= _GEN_395;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_rfSrc2 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_ctrl_rfSrc2 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_ctrl_rfSrc2 <= _GEN_399;
        end
      end else begin
        dataBuffer_3_ctrl_rfSrc2 <= _GEN_399;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_rfWen <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_ctrl_rfWen <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_ctrl_rfWen <= _GEN_403;
        end
      end else begin
        dataBuffer_3_ctrl_rfWen <= _GEN_403;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_rfDest <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_ctrl_rfDest <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_ctrl_rfDest <= _GEN_407;
        end
      end else begin
        dataBuffer_3_ctrl_rfDest <= _GEN_407;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_data_imm <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_7) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_data_imm <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_data_imm <= _GEN_439;
        end
      end else begin
        dataBuffer_3_data_imm <= _GEN_439;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 30:33]
      ringBufferHead <= 2'h0; // @[src/main/scala/utils/PipelineVector.scala 30:33]
    end else if (frontend_io_flushVec[1]) begin // @[src/main/scala/utils/PipelineVector.scala 71:16]
      ringBufferHead <= 2'h0; // @[src/main/scala/utils/PipelineVector.scala 72:24]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      ringBufferHead <= _ringBufferHead_T_1; // @[src/main/scala/utils/PipelineVector.scala 47:24]
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 31:33]
      ringBufferTail <= 2'h0; // @[src/main/scala/utils/PipelineVector.scala 31:33]
    end else if (frontend_io_flushVec[1]) begin // @[src/main/scala/utils/PipelineVector.scala 71:16]
      ringBufferTail <= 2'h0; // @[src/main/scala/utils/PipelineVector.scala 73:24]
    end else if (dequeueFire) begin // @[src/main/scala/utils/PipelineVector.scala 66:22]
      ringBufferTail <= _ringBufferTail_T_1; // @[src/main/scala/utils/PipelineVector.scala 67:24]
    end
    pcOld <= _GEN_1556[31:0]; // @[src/main/scala/nutcore/NutCore.scala 255:{26,26}]
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~someassumeid) begin
          $fwrite(32'h80000002,"Assumption failed\n    at NutCore.scala:132 assume(someAssume)\n"); // @[src/main/scala/nutcore/NutCore.scala 132:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1 & ~_T_19) begin
          $fwrite(32'h80000002,"Assumption failed\n    at NutCore.scala:259 assume(\n"); // @[src/main/scala/nutcore/NutCore.scala 259:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  dataBuffer_0_cf_instr = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  dataBuffer_0_cf_pc = _RAND_1[38:0];
  _RAND_2 = {2{`RANDOM}};
  dataBuffer_0_cf_pnpc = _RAND_2[38:0];
  _RAND_3 = {1{`RANDOM}};
  dataBuffer_0_cf_exceptionVec_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  dataBuffer_0_cf_exceptionVec_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_2 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_3 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_4 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_5 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_6 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_7 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_8 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_9 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_10 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_11 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  dataBuffer_0_cf_brIdx = _RAND_17[3:0];
  _RAND_18 = {1{`RANDOM}};
  dataBuffer_0_ctrl_src1Type = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  dataBuffer_0_ctrl_src2Type = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  dataBuffer_0_ctrl_fuType = _RAND_20[2:0];
  _RAND_21 = {1{`RANDOM}};
  dataBuffer_0_ctrl_fuOpType = _RAND_21[6:0];
  _RAND_22 = {1{`RANDOM}};
  dataBuffer_0_ctrl_rfSrc1 = _RAND_22[4:0];
  _RAND_23 = {1{`RANDOM}};
  dataBuffer_0_ctrl_rfSrc2 = _RAND_23[4:0];
  _RAND_24 = {1{`RANDOM}};
  dataBuffer_0_ctrl_rfWen = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  dataBuffer_0_ctrl_rfDest = _RAND_25[4:0];
  _RAND_26 = {2{`RANDOM}};
  dataBuffer_0_data_imm = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  dataBuffer_1_cf_instr = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  dataBuffer_1_cf_pc = _RAND_28[38:0];
  _RAND_29 = {2{`RANDOM}};
  dataBuffer_1_cf_pnpc = _RAND_29[38:0];
  _RAND_30 = {1{`RANDOM}};
  dataBuffer_1_cf_exceptionVec_1 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  dataBuffer_1_cf_exceptionVec_2 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_0 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_1 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_2 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_3 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_4 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_5 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_6 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_7 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_8 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_9 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_10 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_11 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  dataBuffer_1_cf_brIdx = _RAND_44[3:0];
  _RAND_45 = {1{`RANDOM}};
  dataBuffer_1_ctrl_src1Type = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  dataBuffer_1_ctrl_src2Type = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  dataBuffer_1_ctrl_fuType = _RAND_47[2:0];
  _RAND_48 = {1{`RANDOM}};
  dataBuffer_1_ctrl_fuOpType = _RAND_48[6:0];
  _RAND_49 = {1{`RANDOM}};
  dataBuffer_1_ctrl_rfSrc1 = _RAND_49[4:0];
  _RAND_50 = {1{`RANDOM}};
  dataBuffer_1_ctrl_rfSrc2 = _RAND_50[4:0];
  _RAND_51 = {1{`RANDOM}};
  dataBuffer_1_ctrl_rfWen = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  dataBuffer_1_ctrl_rfDest = _RAND_52[4:0];
  _RAND_53 = {2{`RANDOM}};
  dataBuffer_1_data_imm = _RAND_53[63:0];
  _RAND_54 = {2{`RANDOM}};
  dataBuffer_2_cf_instr = _RAND_54[63:0];
  _RAND_55 = {2{`RANDOM}};
  dataBuffer_2_cf_pc = _RAND_55[38:0];
  _RAND_56 = {2{`RANDOM}};
  dataBuffer_2_cf_pnpc = _RAND_56[38:0];
  _RAND_57 = {1{`RANDOM}};
  dataBuffer_2_cf_exceptionVec_1 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  dataBuffer_2_cf_exceptionVec_2 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_0 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_1 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_2 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_3 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_4 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_5 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_6 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_7 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_8 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_9 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_10 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_11 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  dataBuffer_2_cf_brIdx = _RAND_71[3:0];
  _RAND_72 = {1{`RANDOM}};
  dataBuffer_2_ctrl_src1Type = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  dataBuffer_2_ctrl_src2Type = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  dataBuffer_2_ctrl_fuType = _RAND_74[2:0];
  _RAND_75 = {1{`RANDOM}};
  dataBuffer_2_ctrl_fuOpType = _RAND_75[6:0];
  _RAND_76 = {1{`RANDOM}};
  dataBuffer_2_ctrl_rfSrc1 = _RAND_76[4:0];
  _RAND_77 = {1{`RANDOM}};
  dataBuffer_2_ctrl_rfSrc2 = _RAND_77[4:0];
  _RAND_78 = {1{`RANDOM}};
  dataBuffer_2_ctrl_rfWen = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  dataBuffer_2_ctrl_rfDest = _RAND_79[4:0];
  _RAND_80 = {2{`RANDOM}};
  dataBuffer_2_data_imm = _RAND_80[63:0];
  _RAND_81 = {2{`RANDOM}};
  dataBuffer_3_cf_instr = _RAND_81[63:0];
  _RAND_82 = {2{`RANDOM}};
  dataBuffer_3_cf_pc = _RAND_82[38:0];
  _RAND_83 = {2{`RANDOM}};
  dataBuffer_3_cf_pnpc = _RAND_83[38:0];
  _RAND_84 = {1{`RANDOM}};
  dataBuffer_3_cf_exceptionVec_1 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  dataBuffer_3_cf_exceptionVec_2 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_0 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_1 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_2 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_3 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_4 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_5 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_6 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_7 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_8 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_9 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_10 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_11 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  dataBuffer_3_cf_brIdx = _RAND_98[3:0];
  _RAND_99 = {1{`RANDOM}};
  dataBuffer_3_ctrl_src1Type = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  dataBuffer_3_ctrl_src2Type = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  dataBuffer_3_ctrl_fuType = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  dataBuffer_3_ctrl_fuOpType = _RAND_102[6:0];
  _RAND_103 = {1{`RANDOM}};
  dataBuffer_3_ctrl_rfSrc1 = _RAND_103[4:0];
  _RAND_104 = {1{`RANDOM}};
  dataBuffer_3_ctrl_rfSrc2 = _RAND_104[4:0];
  _RAND_105 = {1{`RANDOM}};
  dataBuffer_3_ctrl_rfWen = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  dataBuffer_3_ctrl_rfDest = _RAND_106[4:0];
  _RAND_107 = {2{`RANDOM}};
  dataBuffer_3_data_imm = _RAND_107[63:0];
  _RAND_108 = {1{`RANDOM}};
  ringBufferHead = _RAND_108[1:0];
  _RAND_109 = {1{`RANDOM}};
  ringBufferTail = _RAND_109[1:0];
  _RAND_110 = {1{`RANDOM}};
  pcOld = _RAND_110[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assume(someassumeid); // @[src/main/scala/nutcore/NutCore.scala 132:9]
    end
    //
    if (_T_1) begin
      assume(_T_19); // @[src/main/scala/nutcore/NutCore.scala 259:13]
    end
  end
endmodule
