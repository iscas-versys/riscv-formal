`define RISCV_FORMAL
`define RISCV_FORMAL_NRET 2
`define RISCV_FORMAL_XLEN 64
`define RISCV_FORMAL_ILEN 32
`define RISCV_FORMAL_RESET_CYCLES 1
`define RISCV_FORMAL_CHECK_CYCLE 20
`define RISCV_FORMAL_CHANNEL_IDX 0
`define RISCV_FORMAL_CHECKER rvfi_insn_check
`define RISCV_FORMAL_INSN_MODEL rvfi_insn_slti
`define RISCV_FORMAL_ALTOPS
`define RISCV_FORMAL_UMODE
`define DEBUGNETS
`define RISCV_FORMAL_COMPRESSED
`include "rvfi_macros.vh"

